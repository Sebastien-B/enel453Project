library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LED_PWM_LUT is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are PWM.

type array_1d is array (0 to 4095) of integer;
constant V2LED_PWM_LUT : array_1d := (

(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(1),
(2),
(4),
(5),
(6),
(8),
(9),
(10),
(12),
(13),
(14),
(16),
(17),
(18),
(19),
(21),
(22),
(23),
(25),
(26),
(27),
(28),
(30),
(31),
(32),
(33),
(35),
(36),
(37),
(38),
(40),
(41),
(42),
(43),
(45),
(46),
(47),
(48),
(49),
(51),
(52),
(53),
(54),
(55),
(57),
(58),
(59),
(60),
(61),
(62),
(64),
(65),
(66),
(67),
(68),
(69),
(71),
(72),
(73),
(74),
(75),
(76),
(77),
(79),
(80),
(81),
(82),
(83),
(84),
(85),
(86),
(88),
(89),
(90),
(91),
(92),
(93),
(94),
(95),
(96),
(97),
(99),
(100),
(101),
(102),
(103),
(104),
(105),
(106),
(107),
(108),
(109),
(110),
(111),
(112),
(113),
(114),
(115),
(117),
(117),
(119),
(120),
(121),
(122),
(123),
(124),
(125),
(126),
(127),
(128),
(129),
(130),
(131),
(132),
(133),
(134),
(135),
(136),
(137),
(138),
(139),
(140),
(141),
(141),
(142),
(143),
(144),
(145),
(146),
(147),
(148),
(149),
(150),
(151),
(152),
(153),
(154),
(155),
(156),
(156),
(157),
(158),
(159),
(160),
(161),
(162),
(163),
(164),
(165),
(166),
(166),
(167),
(168),
(169),
(170),
(171),
(172),
(173),
(173),
(174),
(175),
(176),
(177),
(178),
(179),
(180),
(180),
(181),
(182),
(183),
(184),
(185),
(185),
(186),
(187),
(188),
(189),
(190),
(190),
(191),
(192),
(193),
(194),
(195),
(195),
(196),
(197),
(198),
(199),
(199),
(200),
(201),
(202),
(203),
(203),
(204),
(205),
(206),
(206),
(207),
(208),
(209),
(210),
(210),
(211),
(212),
(213),
(213),
(214),
(215),
(216),
(216),
(217),
(218),
(219),
(219),
(220),
(221),
(222),
(222),
(223),
(224),
(224),
(225),
(226),
(227),
(227),
(228),
(229),
(229),
(230),
(231),
(232),
(232),
(233),
(234),
(234),
(235),
(236),
(236),
(237),
(238),
(239),
(239),
(240),
(240),
(241),
(242),
(243),
(243),
(244),
(245),
(245),
(246),
(247),
(247),
(248),
(248),
(249),
(250),
(250),
(251),
(252),
(252),
(253),
(254),
(254),
(255),
(256),
(256),
(257),
(257),
(258),
(259),
(259),
(260),
(260),
(261),
(262),
(262),
(263),
(263),
(264),
(265),
(265),
(266),
(267),
(267),
(268),
(268),
(269),
(269),
(270),
(271),
(271),
(272),
(272),
(273),
(273),
(274),
(275),
(275),
(276),
(276),
(277),
(277),
(278),
(279),
(279),
(280),
(280),
(281),
(281),
(282),
(282),
(283),
(283),
(284),
(285),
(285),
(286),
(286),
(287),
(287),
(288),
(288),
(289),
(289),
(290),
(290),
(291),
(291),
(292),
(292),
(293),
(293),
(294),
(294),
(295),
(295),
(296),
(296),
(297),
(297),
(298),
(298),
(299),
(299),
(300),
(300),
(301),
(301),
(302),
(302),
(303),
(303),
(304),
(304),
(305),
(305),
(306),
(306),
(307),
(307),
(307),
(308),
(308),
(309),
(309),
(310),
(310),
(311),
(311),
(311),
(312),
(312),
(313),
(313),
(314),
(314),
(315),
(315),
(315),
(316),
(316),
(317),
(317),
(318),
(318),
(319),
(319),
(319),
(320),
(320),
(321),
(321),
(321),
(322),
(322),
(323),
(323),
(323),
(324),
(324),
(325),
(325),
(326),
(326),
(326),
(327),
(327),
(327),
(328),
(328),
(329),
(329),
(329),
(330),
(330),
(331),
(331),
(331),
(332),
(332),
(332),
(333),
(333),
(334),
(334),
(334),
(335),
(335),
(335),
(336),
(336),
(336),
(337),
(337),
(338),
(338),
(338),
(339),
(339),
(339),
(340),
(340),
(340),
(341),
(341),
(341),
(342),
(342),
(343),
(343),
(343),
(343),
(344),
(344),
(344),
(345),
(345),
(346),
(346),
(346),
(347),
(347),
(347),
(347),
(348),
(348),
(348),
(349),
(349),
(349),
(350),
(350),
(350),
(351),
(351),
(351),
(351),
(352),
(352),
(352),
(353),
(353),
(353),
(354),
(354),
(354),
(355),
(355),
(355),
(355),
(356),
(356),
(356),
(357),
(357),
(357),
(358),
(358),
(358),
(358),
(359),
(359),
(359),
(359),
(360),
(360),
(360),
(361),
(361),
(361),
(361),
(362),
(362),
(362),
(362),
(363),
(363),
(363),
(363),
(364),
(364),
(364),
(365),
(365),
(365),
(365),
(366),
(366),
(366),
(366),
(367),
(367),
(367),
(367),
(368),
(368),
(368),
(368),
(369),
(369),
(369),
(369),
(370),
(370),
(370),
(370),
(371),
(371),
(371),
(371),
(372),
(372),
(372),
(372),
(372),
(373),
(373),
(373),
(373),
(374),
(374),
(374),
(374),
(374),
(375),
(375),
(375),
(375),
(376),
(376),
(376),
(376),
(377),
(377),
(377),
(377),
(377),
(378),
(378),
(378),
(378),
(378),
(379),
(379),
(379),
(379),
(379),
(380),
(380),
(380),
(380),
(381),
(381),
(381),
(381),
(381),
(382),
(382),
(382),
(382),
(382),
(382),
(383),
(383),
(383),
(383),
(383),
(384),
(384),
(384),
(384),
(384),
(385),
(385),
(385),
(385),
(385),
(386),
(386),
(386),
(386),
(386),
(386),
(387),
(387),
(387),
(387),
(387),
(388),
(388),
(388),
(388),
(388),
(388),
(389),
(389),
(389),
(389),
(389),
(390),
(390),
(390),
(390),
(390),
(390),
(390),
(391),
(391),
(391),
(391),
(391),
(391),
(392),
(392),
(392),
(392),
(392),
(393),
(393),
(393),
(393),
(393),
(393),
(394),
(394),
(394),
(394),
(394),
(394),
(394),
(394),
(395),
(395),
(395),
(395),
(395),
(395),
(396),
(396),
(396),
(396),
(396),
(396),
(397),
(397),
(397),
(397),
(397),
(397),
(397),
(398),
(398),
(398),
(398),
(398),
(398),
(398),
(398),
(399),
(399),
(399),
(399),
(399),
(399),
(400),
(400),
(400),
(400),
(400),
(400),
(400),
(400),
(401),
(401),
(401),
(401),
(401),
(401),
(401),
(402),
(402),
(402),
(402),
(402),
(402),
(402),
(402),
(403),
(403),
(403),
(403),
(403),
(403),
(403),
(403),
(404),
(404),
(404),
(404),
(404),
(404),
(404),
(405),
(405),
(405),
(405),
(405),
(405),
(405),
(405),
(406),
(406),
(406),
(406),
(406),
(406),
(406),
(406),
(406),
(407),
(407),
(407),
(407),
(407),
(407),
(407),
(407),
(407),
(408),
(408),
(408),
(408),
(408),
(408),
(408),
(408),
(409),
(409),
(409),
(409),
(409),
(409),
(409),
(409),
(409),
(410),
(410),
(410),
(410),
(410),
(410),
(410),
(410),
(410),
(410),
(411),
(411),
(411),
(411),
(411),
(411),
(411),
(411),
(411),
(412),
(412),
(412),
(412),
(412),
(412),
(412),
(412),
(412),
(413),
(413),
(413),
(413),
(413),
(413),
(413),
(413),
(413),
(414),
(414),
(414),
(414),
(414),
(414),
(414),
(414),
(414),
(414),
(414),
(415),
(415),
(415),
(415),
(415),
(415),
(415),
(415),
(415),
(416),
(416),
(416),
(416),
(416),
(416),
(416),
(416),
(416),
(416),
(417),
(417),
(417),
(417),
(417),
(417),
(417),
(417),
(417),
(417),
(418),
(418),
(418),
(418),
(418),
(418),
(418),
(418),
(418),
(418),
(418),
(418),
(419),
(419),
(419),
(419),
(419),
(419),
(419),
(419),
(419),
(419),
(420),
(420),
(420),
(420),
(420),
(420),
(420),
(420),
(420),
(420),
(421),
(421),
(421),
(421),
(421),
(421),
(421),
(421),
(421),
(421),
(422),
(422),
(422),
(422),
(422),
(422),
(422),
(422),
(422),
(422),
(422),
(422),
(423),
(423),
(423),
(423),
(423),
(423),
(423),
(423),
(423),
(423),
(423),
(424),
(424),
(424),
(424),
(424),
(424),
(424),
(424),
(424),
(424),
(425),
(425),
(425),
(425),
(425),
(425),
(425),
(425),
(425),
(425),
(426),
(426),
(426),
(426),
(426),
(426),
(426),
(426),
(426),
(426),
(426),
(426),
(427),
(427),
(427),
(427),
(427),
(427),
(427),
(427),
(427),
(427),
(427),
(428),
(428),
(428),
(428),
(428),
(428),
(428),
(428),
(428),
(428),
(429),
(429),
(429),
(429),
(429),
(429),
(429),
(429),
(429),
(429),
(429),
(430),
(430),
(430),
(430),
(430),
(430),
(430),
(430),
(430),
(430),
(430),
(430),
(431),
(431),
(431),
(431),
(431),
(431),
(431),
(431),
(431),
(431),
(432),
(432),
(432),
(432),
(432),
(432),
(432),
(432),
(432),
(432),
(433),
(433),
(433),
(433),
(433),
(433),
(433),
(433),
(433),
(433),
(434),
(434),
(434),
(434),
(434),
(434),
(434),
(434),
(434),
(434),
(434),
(434),
(435),
(435),
(435),
(435),
(435),
(435),
(435),
(435),
(435),
(435),
(436),
(436),
(436),
(436),
(436),
(436),
(436),
(436),
(436),
(436),
(437),
(437),
(437),
(437),
(437),
(437),
(437),
(437),
(437),
(438),
(438),
(438),
(438),
(438),
(438),
(438),
(438),
(438),
(438),
(438),
(439),
(439),
(439),
(439),
(439),
(439),
(439),
(439),
(439),
(439),
(440),
(440),
(440),
(440),
(440),
(440),
(440),
(440),
(440),
(441),
(441),
(441),
(441),
(441),
(441),
(441),
(441),
(441),
(441),
(442),
(442),
(442),
(442),
(442),
(442),
(442),
(442),
(442),
(442),
(443),
(443),
(443),
(443),
(443),
(443),
(443),
(443),
(443),
(444),
(444),
(444),
(444),
(444),
(444),
(444),
(444),
(444),
(445),
(445),
(445),
(445),
(445),
(445),
(445),
(445),
(445),
(446),
(446),
(446),
(446),
(446),
(446),
(446),
(446),
(446),
(446),
(446),
(447),
(447),
(447),
(447),
(447),
(447),
(447),
(447),
(448),
(448),
(448),
(448),
(448),
(448),
(448),
(448),
(448),
(449),
(449),
(449),
(449),
(449),
(449),
(449),
(449),
(449),
(450),
(450),
(450),
(450),
(450),
(450),
(450),
(450),
(450),
(451),
(451),
(451),
(451),
(451),
(451),
(451),
(451),
(451),
(452),
(452),
(452),
(452),
(452),
(452),
(452),
(452),
(453),
(453),
(453),
(453),
(453),
(453),
(453),
(453),
(454),
(454),
(454),
(454),
(454),
(454),
(454),
(454),
(454),
(454),
(455),
(455),
(455),
(455),
(455),
(455),
(455),
(455),
(456),
(456),
(456),
(456),
(456),
(456),
(456),
(456),
(457),
(457),
(457),
(457),
(457),
(457),
(457),
(457),
(458),
(458),
(458),
(458),
(458),
(458),
(458),
(458),
(458),
(459),
(459),
(459),
(459),
(459),
(459),
(459),
(459),
(460),
(460),
(460),
(460),
(460),
(460),
(460),
(460),
(461),
(461),
(461),
(461),
(461),
(461),
(461),
(461),
(462),
(462),
(462),
(462),
(462),
(462),
(462),
(462),
(463),
(463),
(463),
(463),
(463),
(463),
(463),
(463),
(464),
(464),
(464),
(464),
(464),
(464),
(464),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(465),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(466),
(467),
(467),
(467),
(467),
(467),
(467),
(467),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(468),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(469),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(470),
(471),
(471),
(471),
(471),
(471),
(471),
(471),
(472),
(472),
(472),
(472),
(472),
(472),
(472),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(473),
(474),
(474),
(474),
(474),
(474),
(474),
(474),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(475),
(476),
(476),
(476),
(476),
(476),
(476),
(476),
(477),
(477),
(477),
(477),
(477),
(477),
(477),
(477),
(478),
(478),
(478),
(478),
(478),
(478),
(478),
(478),
(479),
(479),
(479),
(479),
(479),
(479),
(479),
(480),
(480),
(480),
(480),
(480),
(480),
(480),
(480),
(481),
(481),
(481),
(481),
(481),
(481),
(481),
(481),
(482),
(482),
(482),
(482),
(482),
(482),
(482),
(482),
(483),
(483),
(483),
(483),
(483),
(483),
(483),
(484),
(484),
(484),
(484),
(484),
(484),
(484),
(484),
(485),
(485),
(485),
(485),
(485),
(485),
(485),
(485),
(486),
(486),
(486),
(486),
(486),
(486),
(486),
(486),
(487),
(487),
(487),
(487),
(487),
(487),
(487),
(488),
(488),
(488),
(488),
(488),
(488),
(488),
(488),
(489),
(489),
(489),
(489),
(489),
(489),
(489),
(489),
(489),
(490),
(490),
(490),
(490),
(490),
(490),
(490),
(490),
(491),
(491),
(491),
(491),
(491),
(491),
(491),
(491),
(492),
(492),
(492),
(492),
(492),
(492),
(492),
(492),
(493),
(493),
(493),
(493),
(493),
(493),
(493),
(493),
(493),
(494),
(494),
(494),
(494),
(494),
(494),
(494),
(494),
(495),
(495),
(495),
(495),
(495),
(495),
(495),
(495),
(495),
(496),
(496),
(496),
(496),
(496),
(496),
(496),
(496),
(497),
(497),
(497),
(497),
(497),
(497),
(497),
(497),
(497),
(497),
(498),
(498),
(498),
(498),
(498),
(498),
(498),
(498),
(498),
(499),
(499),
(499),
(499),
(499),
(499),
(499),
(499),
(499),
(500),
(500),
(500),
(500),
(500),
(500),
(500),
(500),
(500),
(500),
(501),
(501),
(501),
(501),
(501),
(501),
(501),
(501),
(501),
(501),
(501),
(502),
(502),
(502),
(502),
(502),
(502),
(502),
(502),
(502),
(502),
(503),
(503),
(503),
(503),
(503),
(503),
(503),
(503),
(503),
(503),
(503),
(504),
(504),
(504),
(504),
(504),
(504),
(504),
(504),
(504),
(504),
(504),
(505),
(505),
(505),
(505),
(505),
(505),
(505),
(505),
(505),
(505),
(505),
(505),
(505),
(506),
(506),
(506),
(506),
(506),
(506),
(506),
(506),
(506),
(506),
(506),
(506),
(506),
(507),
(507),
(507),
(507),
(507),
(507),
(507),
(507),
(507),
(507),
(507),
(507),
(507),
(507),
(508),
(508),
(508),
(508),
(508),
(508),
(508),
(508),
(508),
(508),
(508),
(508),
(508),
(508),
(508),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(511),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(510),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(509),
(508),
(508),
(508),
(508),
(508),
(508),
(508),
(508),
(508),
(508),
(508),
(508),
(508),
(507),
(507),
(507),
(507),
(507),
(507),
(507),
(507),
(507),
(507),
(507),
(506),
(506),
(506),
(506),
(506),
(506),
(506),
(506),
(506),
(505),
(505),
(505),
(505),
(505),
(505),
(505),
(505),
(505),
(505),
(504),
(504),
(504),
(504),
(504),
(504),
(504),
(504),
(503),
(503),
(503),
(503),
(503),
(503),
(503),
(502),
(502),
(502),
(502),
(502),
(502),
(502),
(501),
(501),
(501),
(501),
(501),
(501),
(501),
(500),
(500),
(500),
(500),
(500),
(500),
(499),
(499),
(499),
(499),
(499),
(499),
(498),
(498),
(498),
(498),
(498),
(498),
(497),
(497),
(497),
(497),
(497),
(497),
(496),
(496),
(496),
(496),
(496),
(495),
(495),
(495),
(495),
(495),
(494),
(494),
(494),
(494),
(493),
(493),
(493),
(493),
(493),
(492),
(492),
(492),
(492),
(492),
(491),
(491),
(491),
(491),
(490),
(490),
(490),
(490),
(489),
(489),
(489),
(489),
(489),
(488),
(488),
(488),
(488),
(487),
(487),
(487),
(487),
(486),
(486),
(486),
(485),
(485),
(485),
(485),
(485),
(484),
(484),
(484),
(483),
(483),
(483),
(483),
(482),
(482),
(482),
(481),
(481),
(481),
(481),
(480),
(480),
(480),
(479),
(479),
(479),
(478),
(478),
(478),
(478),
(477),
(477),
(477),
(476),
(476),
(476),
(475),
(475),
(475),
(474),
(474),
(474),
(473),
(473),
(473),
(473),
(472),
(472),
(471),
(471),
(471),
(470),
(470),
(470),
(469),
(469),
(469),
(468),
(468),
(468),
(467),
(467),
(466),
(466),
(466),
(465),
(465),
(465),
(464),
(464),
(464),
(463),
(463),
(462),
(462),
(462),
(461),
(461),
(460),
(460),
(460),
(459),
(459),
(458),
(458),
(458),
(457),
(457),
(456),
(456),
(456),
(455),
(455),
(454),
(454),
(453),
(453),
(453),
(452),
(452),
(451),
(451),
(450),
(450),
(450),
(449),
(449),
(448),
(448),
(447),
(447),
(446),
(446),
(445),
(445),
(444),
(444),
(443),
(443),
(442),
(442),
(442),
(441),
(441),
(440),
(440),
(439),
(439),
(438),
(438),
(437),
(437),
(436),
(436),
(435),
(434),
(434),
(434),
(433),
(432),
(432),
(431),
(431),
(430),
(430),
(429),
(429),
(428),
(428),
(427),
(427),
(426),
(426),
(425),
(424),
(424),
(423),
(423),
(422),
(422),
(421),
(420),
(420),
(419),
(419),
(418),
(418),
(417),
(416),
(416),
(415),
(414),
(414),
(413),
(413),
(412),
(411),
(411),
(410),
(410),
(409),
(408),
(408),
(407),
(407),
(406),
(405),
(405),
(404),
(403),
(403),
(402),
(402),
(401),
(400),
(399),
(399),
(398),
(398),
(397),
(396),
(395),
(395),
(394),
(394),
(393),
(392),
(391),
(391),
(390),
(389),
(389),
(388),
(387),
(387),
(386),
(385),
(384),
(384),
(383),
(382),
(382),
(381),
(380),
(379),
(379),
(378),
(377),
(376),
(376),
(375),
(374),
(374),
(373),
(372),
(371),
(370),
(370),
(369),
(368),
(367),
(367),
(366),
(365),
(364),
(363),
(363),
(362),
(361),
(360),
(359),
(359),
(358),
(357),
(356),
(355),
(355),
(354),
(353),
(352),
(351),
(351),
(350),
(349),
(348),
(347),
(346),
(345),
(345),
(344),
(343),
(342),
(341),
(340),
(339),
(339),
(338),
(337),
(336),
(335),
(334),
(333),
(332),
(331),
(331),
(330),
(329),
(328),
(327),
(326),
(325),
(324),
(323),
(322),
(321),
(321),
(320),
(319),
(318),
(317),
(316),
(315),
(314),
(313),
(312),
(311),
(310),
(309),
(308),
(307),
(306),
(305),
(304),
(303),
(302),
(301),
(300),
(299),
(298),
(297),
(296),
(295),
(294),
(293),
(292),
(291),
(290),
(289),
(288),
(287),
(286),
(285),
(284),
(283),
(282),
(281),
(280),
(279),
(278),
(276),
(275),
(274),
(273),
(272),
(271),
(270),
(269),
(268),
(267),
(266),
(264),
(263),
(262),
(261),
(260),
(259),
(258),
(257),
(256),
(254),
(253),
(252),
(251),
(250),
(249),
(247),
(246),
(245),
(244),
(243),
(242),
(240),
(239),
(238),
(237),
(236),
(234),
(233),
(232),
(231),
(230),
(228),
(227),
(226),
(225),
(224),
(222),
(221),
(220),
(219),
(217),
(216),
(215),
(214),
(212),
(211),
(210),
(208),
(207),
(206),
(205),
(203),
(202),
(201),
(200),
(198),
(197),
(196),
(194),
(193),
(192),
(190),
(189),
(188),
(186),
(185),
(184),
(182),
(181),
(180),
(178),
(177),
(176),
(174),
(173),
(171),
(170),
(169),
(167),
(166),
(164),
(163),
(162),
(160),
(159),
(157),
(156),
(155),
(153),
(152),
(150),
(149),
(147),
(146),
(145),
(143),
(142),
(140),
(139),
(137),
(136),
(134),
(133),
(131),
(130),
(128),
(127),
(125),
(124),
(122),
(121),
(119),
(118),
(116),
(115),
(113),
(112),
(110),
(109),
(107),
(105),
(104),
(102),
(101),
(99),
(97),
(96),
(94),
(93),
(91),
(90),
(88),
(86),
(85),
(83),
(82),
(80),
(78),
(77),
(75),
(73),
(72),
(70),
(69),
(67),
(65),
(64),
(62),
(60),
(58),
(57),
(55),
(53),
(52),
(50),
(48),
(47),
(45),
(43),
(42),
(40),
(38),
(36),
(35),
(33),
(31),
(29),
(28),
(26),
(24),
(22),
(21),
(19),
(17),
(15),
(13),
(12),
(10),
(8),
(6),
(4),
(2),
(1),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0),
(0)  -- array index 4095 (voltage = "111111111111" or 4095 mV), distance output 3787 (37.87 cm)
);


end package LED_PWM_LUT;
