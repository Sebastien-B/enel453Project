library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package SEVEN_SEG_PWM_LUT is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are PWM.

type array_1d is array (0 to 4095) of natural;
constant V2SEVEN_SEG_PERIOD_LUT : array_1d := (

--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(488147),
--(487058),
--(485968),
--(484878),
--(483788),
--(482699),
--(481609),
--(480519),
--(479429),
--(478340),
--(477250),
--(476160),
--(475070),
--(473981),
--(472891),
--(471801),
--(470711),
--(469622),
--(468804),
--(467715),
--(466625),
--(465535),
--(464445),
--(463628),
--(462538),
--(461449),
--(460359),
--(459269),
--(458452),
--(457362),
--(456272),
--(455455),
--(454365),
--(453276),
--(452458),
--(451368),
--(450279),
--(449461),
--(448372),
--(447554),
--(446465),
--(445375),
--(444558),
--(443468),
--(442651),
--(441561),
--(440743),
--(439654),
--(438836),
--(437747),
--(436929),
--(435840),
--(435022),
--(433933),
--(433115),
--(432298),
--(431208),
--(430391),
--(429301),
--(428484),
--(427667),
--(426577),
--(425760),
--(424942),
--(423852),
--(423035),
--(422218),
--(421128),
--(420311),
--(419494),
--(418676),
--(417586),
--(416769),
--(415952),
--(415135),
--(414317),
--(413227),
--(412410),
--(411593),
--(410776),
--(409958),
--(409141),
--(408324),
--(407234),
--(406417),
--(405599),
--(404782),
--(403965),
--(403147),
--(402330),
--(401513),
--(400695),
--(399878),
--(399061),
--(398244),
--(397426),
--(396609),
--(395792),
--(394974),
--(394157),
--(393340),
--(392522),
--(391705),
--(390888),
--(390343),
--(389526),
--(388708),
--(387891),
--(387074),
--(386256),
--(385439),
--(384894),
--(384077),
--(383260),
--(382442),
--(381625),
--(381080),
--(380263),
--(379445),
--(378628),
--(378083),
--(377266),
--(376449),
--(375904),
--(375087),
--(374269),
--(373452),
--(372907),
--(372090),
--(371272),
--(370728),
--(369910),
--(369365),
--(368548),
--(367731),
--(367186),
--(366369),
--(365824),
--(365006),
--(364189),
--(363644),
--(362827),
--(362282),
--(361465),
--(360920),
--(360103),
--(359558),
--(358740),
--(358196),
--(357378),
--(356833),
--(356016),
--(355471),
--(354926),
--(354109),
--(353564),
--(352747),
--(352202),
--(351385),
--(350840),
--(350295),
--(349478),
--(348933),
--(348388),
--(347571),
--(347026),
--(346481),
--(345663),
--(345119),
--(344574),
--(343756),
--(343212),
--(342667),
--(342122),
--(341305),
--(340760),
--(340215),
--(339670),
--(338853),
--(338308),
--(337763),
--(337218),
--(336673),
--(335856),
--(335311),
--(334766),
--(334221),
--(333676),
--(333131),
--(332314),
--(331769),
--(331224),
--(330680),
--(330135),
--(329590),
--(329045),
--(328500),
--(327683),
--(327138),
--(326593),
--(326048),
--(325503),
--(324958),
--(324414),
--(323869),
--(323324),
--(322779),
--(322234),
--(321689),
--(321144),
--(320599),
--(320055),
--(319510),
--(318965),
--(318420),
--(317875),
--(317330),
--(316785),
--(316240),
--(315968),
--(315423),
--(314878),
--(314333),
--(313789),
--(313244),
--(312699),
--(312154),
--(311609),
--(311337),
--(310792),
--(310247),
--(309702),
--(309157),
--(308612),
--(308067),
--(307795),
--(307250),
--(306705),
--(306160),
--(305615),
--(305343),
--(304798),
--(304253),
--(303708),
--(303436),
--(302891),
--(302346),
--(301801),
--(301529),
--(300984),
--(300439),
--(299894),
--(299622),
--(299077),
--(298532),
--(298260),
--(297715),
--(297170),
--(296898),
--(296353),
--(295808),
--(295535),
--(294990),
--(294446),
--(294173),
--(293628),
--(293356),
--(292811),
--(292266),
--(291994),
--(291449),
--(290904),
--(290632),
--(290087),
--(289814),
--(289269),
--(288997),
--(288452),
--(287907),
--(287635),
--(287090),
--(286817),
--(286273),
--(286000),
--(285455),
--(285183),
--(284638),
--(284365),
--(283821),
--(283548),
--(283003),
--(282731),
--(282186),
--(281914),
--(281369),
--(281096),
--(280551),
--(280279),
--(280007),
--(279462),
--(279189),
--(278644),
--(278372),
--(277827),
--(277555),
--(277282),
--(276737),
--(276465),
--(275920),
--(275648),
--(275375),
--(274830),
--(274558),
--(274013),
--(273741),
--(273468),
--(272923),
--(272651),
--(272378),
--(271833),
--(271561),
--(271289),
--(270744),
--(270471),
--(270199),
--(269654),
--(269382),
--(269109),
--(268564),
--(268292),
--(268019),
--(267747),
--(267202),
--(266930),
--(266657),
--(266112),
--(265840),
--(265567),
--(265295),
--(264750),
--(264478),
--(264205),
--(263933),
--(263388),
--(263116),
--(262843),
--(262571),
--(262298),
--(261753),
--(261481),
--(261208),
--(260936),
--(260664),
--(260119),
--(259846),
--(259574),
--(259301),
--(259029),
--(258484),
--(258212),
--(257939),
--(257667),
--(257394),
--(257122),
--(256577),
--(256305),
--(256032),
--(255760),
--(255487),
--(255215),
--(254942),
--(254670),
--(254125),
--(253853),
--(253580),
--(253308),
--(253035),
--(252763),
--(252491),
--(252218),
--(251946),
--(251673),
--(251128),
--(250856),
--(250583),
--(250311),
--(250039),
--(249766),
--(249494),
--(249221),
--(248949),
--(248676),
--(248404),
--(248132),
--(247859),
--(247587),
--(247314),
--(247042),
--(246769),
--(246497),
--(246225),
--(245952),
--(245680),
--(245135),
--(244862),
--(244590),
--(244317),
--(244045),
--(243773),
--(243500),
--(243228),
--(243228),
--(242955),
--(242683),
--(242410),
--(242138),
--(241866),
--(241593),
--(241321),
--(241048),
--(240776),
--(240503),
--(240231),
--(239958),
--(239686),
--(239414),
--(239141),
--(238869),
--(238596),
--(238324),
--(238051),
--(237779),
--(237507),
--(237234),
--(237234),
--(236962),
--(236689),
--(236417),
--(236144),
--(235872),
--(235600),
--(235327),
--(235055),
--(234782),
--(234510),
--(234510),
--(234237),
--(233965),
--(233692),
--(233420),
--(233148),
--(232875),
--(232603),
--(232603),
--(232330),
--(232058),
--(231785),
--(231513),
--(231241),
--(230968),
--(230696),
--(230696),
--(230423),
--(230151),
--(229878),
--(229606),
--(229334),
--(229061),
--(229061),
--(228789),
--(228516),
--(228244),
--(227971),
--(227699),
--(227699),
--(227426),
--(227154),
--(226882),
--(226609),
--(226609),
--(226337),
--(226064),
--(225792),
--(225519),
--(225247),
--(225247),
--(224975),
--(224702),
--(224430),
--(224157),
--(224157),
--(223885),
--(223612),
--(223340),
--(223067),
--(223067),
--(222795),
--(222523),
--(222250),
--(222250),
--(221978),
--(221705),
--(221433),
--(221160),
--(221160),
--(220888),
--(220616),
--(220343),
--(220343),
--(220071),
--(219798),
--(219526),
--(219253),
--(219253),
--(218981),
--(218709),
--(218436),
--(218436),
--(218164),
--(217891),
--(217619),
--(217619),
--(217346),
--(217074),
--(216801),
--(216801),
--(216529),
--(216257),
--(215984),
--(215984),
--(215712),
--(215439),
--(215439),
--(215167),
--(214894),
--(214622),
--(214622),
--(214350),
--(214077),
--(213805),
--(213805),
--(213532),
--(213260),
--(212987),
--(212987),
--(212715),
--(212443),
--(212443),
--(212170),
--(211898),
--(211625),
--(211625),
--(211353),
--(211080),
--(211080),
--(210808),
--(210535),
--(210263),
--(210263),
--(209991),
--(209718),
--(209718),
--(209446),
--(209173),
--(209173),
--(208901),
--(208628),
--(208356),
--(208356),
--(208084),
--(207811),
--(207811),
--(207539),
--(207266),
--(207266),
--(206994),
--(206721),
--(206449),
--(206449),
--(206176),
--(205904),
--(205904),
--(205632),
--(205359),
--(205359),
--(205087),
--(204814),
--(204814),
--(204542),
--(204269),
--(204269),
--(203997),
--(203725),
--(203452),
--(203452),
--(203180),
--(202907),
--(202907),
--(202635),
--(202362),
--(202362),
--(202090),
--(201818),
--(201818),
--(201545),
--(201273),
--(201273),
--(201000),
--(200728),
--(200728),
--(200455),
--(200183),
--(200183),
--(199910),
--(199638),
--(199638),
--(199366),
--(199093),
--(199093),
--(198821),
--(198548),
--(198548),
--(198276),
--(198003),
--(198003),
--(197731),
--(197459),
--(197459),
--(197186),
--(196914),
--(196914),
--(196641),
--(196369),
--(196096),
--(196096),
--(195824),
--(195552),
--(195552),
--(195279),
--(195007),
--(195007),
--(194734),
--(194462),
--(194462),
--(194189),
--(193917),
--(193917),
--(193644),
--(193372),
--(193372),
--(193100),
--(192827),
--(192827),
--(192555),
--(192282),
--(192282),
--(192010),
--(191737),
--(191737),
--(191465),
--(191193),
--(191193),
--(190920),
--(190648),
--(190648),
--(190375),
--(190103),
--(190103),
--(189830),
--(189558),
--(189558),
--(189285),
--(189013),
--(189013),
--(188741),
--(188468),
--(188468),
--(188196),
--(187923),
--(187923),
--(187651),
--(187378),
--(187378),
--(187106),
--(186834),
--(186834),
--(186561),
--(186289),
--(186289),
--(186016),
--(185744),
--(185744),
--(185471),
--(185199),
--(185199),
--(184927),
--(184654),
--(184654),
--(184382),
--(184109),
--(184109),
--(183837),
--(183564),
--(183564),
--(183292),
--(183019),
--(183019),
--(182747),
--(182475),
--(182202),
--(182202),
--(181930),
--(181657),
--(181657),
--(181385),
--(181112),
--(181112),
--(180840),
--(180568),
--(180568),
--(180295),
--(180023),
--(180023),
--(179750),
--(179478),
--(179478),
--(179205),
--(178933),
--(178661),
--(178661),
--(178388),
--(178116),
--(178116),
--(177843),
--(177571),
--(177571),
--(177298),
--(177026),
--(177026),
--(176753),
--(176481),
--(176209),
--(176209),
--(175936),
--(175664),
--(175664),
--(175391),
--(175119),
--(175119),
--(174846),
--(174574),
--(174302),
--(174302),
--(174029),
--(173757),
--(173757),
--(173484),
--(173212),
--(172939),
--(172939),
--(172667),
--(172394),
--(172394),
--(172122),
--(171850),
--(171850),
--(171577),
--(171305),
--(171032),
--(171032),
--(170760),
--(170487),
--(170215),
--(170215),
--(169943),
--(169670),
--(169670),
--(169398),
--(169125),
--(168853),
--(168853),
--(168580),
--(168308),
--(168308),
--(168036),
--(167763),
--(167491),
--(167491),
--(167218),
--(166946),
--(166673),
--(166673),
--(166401),
--(166128),
--(166128),
--(165856),
--(165584),
--(165311),
--(165311),
--(165039),
--(164766),
--(164494),
--(164494),
--(164221),
--(163949),
--(163677),
--(163677),
--(163404),
--(163132),
--(162859),
--(162859),
--(162587),
--(162314),
--(162042),
--(162042),
--(161770),
--(161497),
--(161225),
--(161225),
--(160952),
--(160680),
--(160407),
--(160407),
--(160135),
--(159862),
--(159590),
--(159590),
--(159318),
--(159045),
--(158773),
--(158773),
--(158500),
--(158228),
--(157955),
--(157683),
--(157683),
--(157411),
--(157138),
--(156866),
--(156866),
--(156593),
--(156321),
--(156048),
--(155776),
--(155776),
--(155503),
--(155231),
--(154959),
--(154959),
--(154686),
--(154414),
--(154141),
--(153869),
--(153869),
--(153596),
--(153324),
--(153052),
--(152779),
--(152779),
--(152507),
--(152234),
--(151962),
--(151962),
--(151689),
--(151417),
--(151145),
--(150872),
--(150872),
--(150600),
--(150327),
--(150055),
--(149782),
--(149782),
--(149510),
--(149237),
--(148965),
--(148693),
--(148693),
--(148420),
--(148148),
--(147875),
--(147603),
--(147330),
--(147330),
--(147058),
--(146786),
--(146513),
--(146241),
--(146241),
--(145968),
--(145696),
--(145423),
--(145151),
--(144879),
--(144879),
--(144606),
--(144334),
--(144061),
--(143789),
--(143516),
--(143516),
--(143244),
--(142971),
--(142699),
--(142427),
--(142154),
--(142154),
--(141882),
--(141609),
--(141337),
--(141064),
--(140792),
--(140792),
--(140520),
--(140247),
--(139975),
--(139702),
--(139430),
--(139430),
--(139157),
--(138885),
--(138612),
--(138340),
--(138068),
--(137795),
--(137795),
--(137523),
--(137250),
--(136978),
--(136705),
--(136433),
--(136161),
--(136161),
--(135888),
--(135616),
--(135343),
--(135071),
--(134798),
--(134526),
--(134526),
--(134254),
--(133981),
--(133709),
--(133436),
--(133164),
--(132891),
--(132619),
--(132619),
--(132346),
--(132074),
--(131802),
--(131529),
--(131257),
--(130984),
--(130712),
--(130712),
--(130439),
--(130167),
--(129895),
--(129622),
--(129350),
--(129077),
--(128805),
--(128805),
--(128532),
--(128260),
--(127987),
--(127715),
--(127443),
--(127170),
--(126898),
--(126625),
--(126625),
--(126353),
--(126080),
--(125808),
--(125536),
--(125263),
--(124991),
--(124718),
--(124446),
--(124446),
--(124173),
--(123901),
--(123629),
--(123356),
--(123084),
--(122811),
--(122539),
--(122266),
--(121994),
--(121721),
--(121721),
--(121449),
--(121177),
--(120904),
--(120632),
--(120359),
--(120087),
--(119814),
--(119542),
--(119270),
--(118997),
--(118997),
--(118725),
--(118452),
--(118180),
--(117907),
--(117635),
--(117363),
--(117090),
--(116818),
--(116545),
--(116273),
--(116000),
--(116000),
--(115728),
--(115455),
--(115183),
--(114911),
--(114638),
--(114366),
--(114093),
--(113821),
--(113548),
--(113276),
--(113004),
--(112731),
--(112731),
--(112459),
--(112186),
--(111914),
--(111641),
--(111369),
--(111096),
--(110824),
--(110552),
--(110279),
--(110007),
--(109734),
--(109462),
--(109189),
--(108917),
--(108917),
--(108645),
--(108372),
--(108100),
--(107827),
--(107555),
--(107282),
--(107010),
--(106738),
--(106465),
--(106193),
--(105920),
--(105648),
--(105375),
--(105103),
--(104830),
--(104830),
--(104558),
--(104286),
--(104013),
--(103741),
--(103468),
--(103196),
--(102923),
--(102651),
--(102379),
--(102106),
--(101834),
--(101561),
--(101289),
--(101016),
--(100744),
--(100472),
--(100199),
--(100199),
--(99927),
--(99654),
--(99382),
--(99109),
--(98837),
--(98564),
--(98292),
--(98020),
--(97747),
--(97475),
--(97202),
--(96930),
--(96657),
--(96385),
--(96113),
--(95840),
--(95568),
--(95295),
--(95295),
--(95023),
--(94750),
--(94478),
--(94205),
--(93933),
--(93661),
--(93388),
--(93116),
--(92843),
--(92571),
--(92298),
--(92026),
--(91754),
--(91481),
--(91209),
--(90936),
--(90664),
--(90391),
--(90119),
--(90119),
--(89847),
--(89574),
--(89302),
--(89029),
--(88757),
--(88484),
--(88212),
--(87939),
--(87667),
--(87395),
--(87122),
--(86850),
--(86577),
--(86305),
--(86032),
--(85760),
--(85488),
--(85488),
--(85215),
--(84943),
--(84670),
--(84398),
--(84125),
--(83853),
--(83581),
--(83308),
--(83036),
--(82763),
--(82491),
--(82218),
--(81946),
--(81673),
--(81401),
--(81129),
--(80856),
--(80856),
--(80584),
--(80311),
--(80039),
--(79766),
--(79494),
--(79222),
--(78949),
--(78677),
--(78404),
--(78132),
--(77859),
--(77587),
--(77314),
--(77042),
--(77042),
--(76770),
--(76497),
--(76225),
--(75952),
--(75680),
--(75407),
--(75135),
--(74863),
--(74590),
--(74318),
--(74045),
--(73773),
--(73773),
--(73500),
--(73228),
--(72956),
--(72683),
--(72411),
--(72138),
--(71866),
--(71593),
--(71321),
--(71048),
--(70776),
--(70776),
--(70504),
--(70231),
--(69959),
--(69686),
--(69414),
--(69141),
--(68869),
--(68597),
--(68324),
--(68052),
--(68052),
--(67779),
--(67507),
--(67234),
--(66962),
--(66690),
--(66417),
--(66145),
--(65872),
--(65600),
--(65600),
--(65327),
--(65055),
--(64782),
--(64510),
--(64238),
--(63965),
--(63693),
--(63693),
--(63420),
--(63148),
--(62875),
--(62603),
--(62331),
--(62058),
--(61786),
--(61786),
--(61513),
--(61241),
--(60968),
--(60696),
--(60423),
--(60151),
--(59879),
--(59879),
--(59606),
--(59334),
--(59061),
--(58789),
--(58516),
--(58244),
--(58244),
--(57972),
--(57699),
--(57427),
--(57154),
--(56882),
--(56882),
--(56609),
--(56337),
--(56065),
--(55792),
--(55520),
--(55520),
--(55247),
--(54975),
--(54702),
--(54430),
--(54157),
--(54157),
--(53885),
--(53613),
--(53340),
--(53068),
--(53068),
--(52795),
--(52523),
--(52250),
--(51978),
--(51706),
--(51706),
--(51433),
--(51161),
--(50888),
--(50888),
--(50616),
--(50343),
--(50071),
--(49799),
--(49799),
--(49526),
--(49254),
--(48981),
--(48709),
--(48709),
--(48436),
--(48164),
--(47891),
--(47891),
--(47619),
--(47347),
--(47074),
--(47074),
--(46802),
--(46529),
--(46257),
--(46257),
--(45984),
--(45712),
--(45440),
--(45440),
--(45167),
--(44895),
--(44622),
--(44622),
--(44350),
--(44077),
--(44077),
--(43805),
--(43532),
--(43260),
--(43260),
--(42988),
--(42715),
--(42715),
--(42443),
--(42170),
--(42170),
--(41898),
--(41625),
--(41353),
--(41353),
--(41081),
--(40808),
--(40808),
--(40536),
--(40263),
--(40263),
--(39991),
--(39718),
--(39718),
--(39446),
--(39446),
--(39174),
--(38901),
--(38901),
--(38629),
--(38356),
--(38356),
--(38084),
--(37811),
--(37811),
--(37539),
--(37539),
--(37266),
--(36994),
--(36994),
--(36722),
--(36722),
--(36449),
--(36177),
--(36177),
--(35904),
--(35904),
--(35632),
--(35359),
--(35359),
--(35087),
--(35087),
--(34815),
--(34815),
--(34542),
--(34270),
--(34270),
--(33997),
--(33997),
--(33725),
--(33725),
--(33452),
--(33452),
--(33180),
--(33180),
--(32908),
--(32908),
--(32635),
--(32635),
--(32363),
--(32090),
--(32090),
--(31818),
--(31818),
--(31818),
--(31545),
--(31545),
--(31273),
--(31273),
--(31000),
--(31000),
--(30728),
--(30728),
--(30456),
--(30456),
--(30183),
--(30183),
--(30183),
--(29911),
--(29911),
--(29638),
--(29638),
--(29366),
--(29366),
--(29366),
--(29093),
--(29093),
--(28821),
--(28821),
--(28821),
--(28549),
--(28549),
--(28276),
--(28276),
--(28276),
--(28004),
--(28004),
--(28004),
--(27731),
--(27731),
--(27731),
--(27459),
--(27459),
--(27459),
--(27186),
--(27186),
--(27186),
--(26914),
--(26914),
--(26914),
--(26641),
--(26641),
--(26641),
--(26641),
--(26369),
--(26369),
--(26369),
--(26369),
--(26097),
--(26097),
--(26097),
--(26097),
--(25824),
--(25824),
--(25824),
--(25824),
--(25552),
--(25552),
--(25552),
--(25552),
--(25552),
--(25279),
--(25279),
--(25279),
--(25279),
--(25279),
--(25007),
--(25007),
--(25007),
--(25007),
--(25007),
--(25007),
--(25007),
--(24734),
--(24734),
--(24734),
--(24734),
--(24734),
--(24734),
--(24734),
--(24734),
--(24734),
--(24734),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24462),
--(24734),
--(24734),
--(24734),
--(24734),
--(24734),
--(24734),
--(24734),
--(24734),
--(24734),
--(25007),
--(25007),
--(25007),
--(25007),
--(25007),
--(25007),
--(25279),
--(25279),
--(25279),
--(25279),
--(25279),
--(25552),
--(25552),
--(25552),
--(25552),
--(25552),
--(25824),
--(25824),
--(25824),
--(25824),
--(26097),
--(26097),
--(26097),
--(26369),
--(26369),
--(26369),
--(26369),
--(26641),
--(26641),
--(26641),
--(26914),
--(26914),
--(26914),
--(27186),
--(27186),
--(27459),
--(27459),
--(27459),
--(27731),
--(27731),
--(28004),
--(28004),
--(28004),
--(28276),
--(28276),
--(28549),
--(28549),
--(28821),
--(28821),
--(29093),
--(29093),
--(29366),
--(29366),
--(29638),
--(29638),
--(29911),
--(29911),
--(30183),
--(30183),
--(30456),
--(30456),
--(30728),
--(31000),
--(31000),
--(31273),
--(31273),
--(31545),
--(31818),
--(31818),
--(32090),
--(32090),
--(32363),
--(32635),
--(32635),
--(32908),
--(33180),
--(33180),
--(33452),
--(33725),
--(33997),
--(33997),
--(34270),
--(34542),
--(34542),
--(34815),
--(35087),
--(35359),
--(35632),
--(35632),
--(35904),
--(36177),
--(36449),
--(36722),
--(36722),
--(36994),
--(37266),
--(37539),
--(37811),
--(38084),
--(38356),
--(38629),
--(38629),
--(38901),
--(39174),
--(39446),
--(39718),
--(39991),
--(40263),
--(40536),
--(40808),
--(41081),
--(41353),
--(41625),
--(41898),
--(42170),
--(42443),
--(42715),
--(42988),
--(43260),
--(43532),
--(43805),
--(44077),
--(44350),
--(44895),
--(45167),
--(45440),
--(45712),
--(45984),
--(46257),
--(46529),
--(47074),
--(47347),
--(47619),
--(47891),
--(48164),
--(48709),
--(48981),
--(49254),
--(49526),
--(50071),
--(50343),
--(50616),
--(50888),
--(51433),
--(51706),
--(51978),
--(52523),
--(52795),
--(53068),
--(53613),
--(53885),
--(54157),
--(54702),
--(54975),
--(55520),
--(55792),
--(56337),
--(56609),
--(56882),
--(57427),
--(57699),
--(58244),
--(58516),
--(59061),
--(59334),
--(59879),
--(60151),
--(60696),
--(61241),
--(61513),
--(62058),
--(62331),
--(62875),
--(63420),
--(63693),
--(64238),
--(64510),
--(65055),
--(65600),
--(65872),
--(66417),
--(66962),
--(67507),
--(67779),
--(68324),
--(68869),
--(69414),
--(69686),
--(70231),
--(70776),
--(71321),
--(71593),
--(72138),
--(72683),
--(73228),
--(73773),
--(74318),
--(74863),
--(75135),
--(75680),
--(76225),
--(76770),
--(77314),
--(77859),
--(78404),
--(78949),
--(79494),
--(80039),
--(80584),
--(81129),
--(81673),
--(82218),
--(82763),
--(83308),
--(83853),
--(84670),
--(85215),
--(85760),
--(86305),
--(86850),
--(87395),
--(87939),
--(88757),
--(89302),
--(89847),
--(90391),
--(90936),
--(91754),
--(92298),
--(92843),
--(93388),
--(94205),
--(94750),
--(95295),
--(96113),
--(96657),
--(97202),
--(98020),
--(98564),
--(99382),
--(99927),
--(100472),
--(101289),
--(101834),
--(102651),
--(103196),
--(104013),
--(104558),
--(105375),
--(105920),
--(106738),
--(107282),
--(108100),
--(108917),
--(109462),
--(110279),
--(110824),
--(111641),
--(112459),
--(113004),
--(113821),
--(114638),
--(115183),
--(116000),
--(116818),
--(117635),
--(118180),
--(118997),
--(119814),
--(120632),
--(121177),
--(121994),
--(122811),
--(123629),
--(124446),
--(125263),
--(126080),
--(126898),
--(127443),
--(128260),
--(129077),
--(129895),
--(130712),
--(131529),
--(132346),
--(133164),
--(133981),
--(134798),
--(135888),
--(136705),
--(137523),
--(138340),
--(139157),
--(139975),
--(140792),
--(141609),
--(142699),
--(143516),
--(144334),
--(145151),
--(145968),
--(147058),
--(147875),
--(148693),
--(149782),
--(150600),
--(151417),
--(152507),
--(153324),
--(154141),
--(155231),
--(156048),
--(157138),
--(157955),
--(158773),
--(159862),
--(160680),
--(161770),
--(162587),
--(163677),
--(164766),
--(165584),
--(166673),
--(167491),
--(168580),
--(169670),
--(170487),
--(171577),
--(172667),
--(173484),
--(174574),
--(175664),
--(176481),
--(177571),
--(178661),
--(179750),
--(180840),
--(181657),
--(182747),
--(183837),
--(184927),
--(186016),
--(187106),
--(188196),
--(189285),
--(190103),
--(191193),
--(192282),
--(193372),
--(194462),
--(195552),
--(196914),
--(198003),
--(199093),
--(200183),
--(201273),
--(202362),
--(203452),
--(204542),
--(205904),
--(206994),
--(208084),
--(209173),
--(210263),
--(211625),
--(212715),
--(213805),
--(215167),
--(216257),
--(217346),
--(218709),
--(219798),
--(221160),
--(222250),
--(223340),
--(224702),
--(225792),
--(227154),
--(228244),
--(229606),
--(230696),
--(232058),
--(233420),
--(234510),
--(235872),
--(236962),
--(238324),
--(239686),
--(240776),
--(242138),
--(243500),
--(244862),
--(245952),
--(247314),
--(248676),
--(250039),
--(251401),
--(252763),
--(253853),
--(255215),
--(256577),
--(257939),
--(259301),
--(260664),
--(262026),
--(263388),
--(264750),
--(266112),
--(267474),
--(268837),
--(270199),
--(271561),
--(273196),
--(274558),
--(275920),
--(277282),
--(278644),
--(280279),
--(281641),
--(283003),
--(284365),
--(286000),
--(287362),
--(288724),
--(290359),
--(291721),
--(293356),
--(294718),
--(296080),
--(297715),
--(299077),
--(300712),
--(302074),
--(303708),
--(305071),
--(306705),
--(308340),
--(309702),
--(311337),
--(312971),
--(314333),
--(315968),
--(317603),
--(318965),
--(320599),
--(322234),
--(323869),
--(325503),
--(326865),
--(328500),
--(330135),
--(331769),
--(333404),
--(335038),
--(336673),
--(338308),
--(339942),
--(341577),
--(343212),
--(344846),
--(346481),
--(348115),
--(349750),
--(351657),
--(353292),
--(354926),
--(356561),
--(358196),
--(360103),
--(361737),
--(363372),
--(365279),
--(366913),
--(368548),
--(370455),
--(372090),
--(373724),
--(375631),
--(377266),
--(379173),
--(380808),
--(382715),
--(384349),
--(386256),
--(388163),
--(389798),
--(391705),
--(393612),
--(395247),
--(397154),
--(399061),
--(400695),
--(402603),
--(404510),
--(406417),
--(408324),
--(410231),
--(411865),
--(413772),
--(415679),
--(417586),
--(419494),
--(421401),
--(423308),
--(425215),
--(427122),
--(429029),
--(431208),
--(433115),
--(435022),
--(436929),
--(438836),
--(441016),
--(442923),
--(444830),
--(446737),
--(448917),
--(450824),
--(452731),
--(454910),
--(456817),
--(458997),
--(460904),
--(463083),
--(464990),
--(467170),
--(469077),
--(471256),
--(473163),
--(475343),
--(477522),
--(479429),
--(481609),
--(483788),
--(485695),
--(487875),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237),
--(489237)  -- array index 4095 (voltage = "111111111111" or 4095 mV), distance output 3787 (37.87 cm)

(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	162	)	,
(	162	)	,
(	161	)	,
(	161	)	,
(	161	)	,
(	160	)	,
(	160	)	,
(	159	)	,
(	159	)	,
(	159	)	,
(	158	)	,
(	158	)	,
(	157	)	,
(	157	)	,
(	157	)	,
(	156	)	,
(	156	)	,
(	156	)	,
(	155	)	,
(	155	)	,
(	154	)	,
(	154	)	,
(	154	)	,
(	153	)	,
(	153	)	,
(	153	)	,
(	152	)	,
(	152	)	,
(	151	)	,
(	151	)	,
(	151	)	,
(	150	)	,
(	150	)	,
(	150	)	,
(	149	)	,
(	149	)	,
(	148	)	,
(	148	)	,
(	148	)	,
(	147	)	,
(	147	)	,
(	147	)	,
(	146	)	,
(	146	)	,
(	146	)	,
(	145	)	,
(	145	)	,
(	145	)	,
(	144	)	,
(	144	)	,
(	143	)	,
(	143	)	,
(	143	)	,
(	142	)	,
(	142	)	,
(	142	)	,
(	141	)	,
(	141	)	,
(	141	)	,
(	140	)	,
(	140	)	,
(	140	)	,
(	139	)	,
(	139	)	,
(	139	)	,
(	138	)	,
(	138	)	,
(	138	)	,
(	137	)	,
(	137	)	,
(	137	)	,
(	136	)	,
(	136	)	,
(	136	)	,
(	135	)	,
(	135	)	,
(	135	)	,
(	134	)	,
(	134	)	,
(	134	)	,
(	133	)	,
(	133	)	,
(	133	)	,
(	132	)	,
(	132	)	,
(	132	)	,
(	132	)	,
(	131	)	,
(	131	)	,
(	131	)	,
(	130	)	,
(	130	)	,
(	130	)	,
(	129	)	,
(	129	)	,
(	129	)	,
(	128	)	,
(	128	)	,
(	128	)	,
(	127	)	,
(	127	)	,
(	127	)	,
(	127	)	,
(	126	)	,
(	126	)	,
(	126	)	,
(	125	)	,
(	125	)	,
(	125	)	,
(	124	)	,
(	124	)	,
(	124	)	,
(	124	)	,
(	123	)	,
(	123	)	,
(	123	)	,
(	122	)	,
(	122	)	,
(	122	)	,
(	121	)	,
(	121	)	,
(	121	)	,
(	121	)	,
(	120	)	,
(	120	)	,
(	120	)	,
(	119	)	,
(	119	)	,
(	119	)	,
(	119	)	,
(	118	)	,
(	118	)	,
(	118	)	,
(	118	)	,
(	117	)	,
(	117	)	,
(	117	)	,
(	116	)	,
(	116	)	,
(	116	)	,
(	116	)	,
(	115	)	,
(	115	)	,
(	115	)	,
(	114	)	,
(	114	)	,
(	114	)	,
(	114	)	,
(	113	)	,
(	113	)	,
(	113	)	,
(	113	)	,
(	112	)	,
(	112	)	,
(	112	)	,
(	112	)	,
(	111	)	,
(	111	)	,
(	111	)	,
(	111	)	,
(	110	)	,
(	110	)	,
(	110	)	,
(	109	)	,
(	109	)	,
(	109	)	,
(	109	)	,
(	108	)	,
(	108	)	,
(	108	)	,
(	108	)	,
(	107	)	,
(	107	)	,
(	107	)	,
(	107	)	,
(	106	)	,
(	106	)	,
(	106	)	,
(	106	)	,
(	105	)	,
(	105	)	,
(	105	)	,
(	105	)	,
(	105	)	,
(	104	)	,
(	104	)	,
(	104	)	,
(	104	)	,
(	103	)	,
(	103	)	,
(	103	)	,
(	103	)	,
(	102	)	,
(	102	)	,
(	102	)	,
(	102	)	,
(	101	)	,
(	101	)	,
(	101	)	,
(	101	)	,
(	100	)	,
(	100	)	,
(	100	)	,
(	100	)	,
(	100	)	,
(	99	)	,
(	99	)	,
(	99	)	,
(	99	)	,
(	98	)	,
(	98	)	,
(	98	)	,
(	98	)	,
(	98	)	,
(	97	)	,
(	97	)	,
(	97	)	,
(	97	)	,
(	96	)	,
(	96	)	,
(	96	)	,
(	96	)	,
(	96	)	,
(	95	)	,
(	95	)	,
(	95	)	,
(	95	)	,
(	95	)	,
(	94	)	,
(	94	)	,
(	94	)	,
(	94	)	,
(	93	)	,
(	93	)	,
(	93	)	,
(	93	)	,
(	93	)	,
(	92	)	,
(	92	)	,
(	92	)	,
(	92	)	,
(	92	)	,
(	91	)	,
(	91	)	,
(	91	)	,
(	91	)	,
(	91	)	,
(	90	)	,
(	90	)	,
(	90	)	,
(	90	)	,
(	90	)	,
(	89	)	,
(	89	)	,
(	89	)	,
(	89	)	,
(	89	)	,
(	88	)	,
(	88	)	,
(	88	)	,
(	88	)	,
(	88	)	,
(	87	)	,
(	87	)	,
(	87	)	,
(	87	)	,
(	87	)	,
(	87	)	,
(	86	)	,
(	86	)	,
(	86	)	,
(	86	)	,
(	86	)	,
(	85	)	,
(	85	)	,
(	85	)	,
(	85	)	,
(	85	)	,
(	85	)	,
(	84	)	,
(	84	)	,
(	84	)	,
(	84	)	,
(	84	)	,
(	83	)	,
(	83	)	,
(	83	)	,
(	83	)	,
(	83	)	,
(	83	)	,
(	82	)	,
(	82	)	,
(	82	)	,
(	82	)	,
(	82	)	,
(	82	)	,
(	81	)	,
(	81	)	,
(	81	)	,
(	81	)	,
(	81	)	,
(	81	)	,
(	80	)	,
(	80	)	,
(	80	)	,
(	80	)	,
(	80	)	,
(	80	)	,
(	79	)	,
(	79	)	,
(	79	)	,
(	79	)	,
(	79	)	,
(	79	)	,
(	78	)	,
(	78	)	,
(	78	)	,
(	78	)	,
(	78	)	,
(	78	)	,
(	77	)	,
(	77	)	,
(	77	)	,
(	77	)	,
(	77	)	,
(	77	)	,
(	76	)	,
(	76	)	,
(	76	)	,
(	76	)	,
(	76	)	,
(	76	)	,
(	76	)	,
(	75	)	,
(	75	)	,
(	75	)	,
(	75	)	,
(	75	)	,
(	75	)	,
(	74	)	,
(	74	)	,
(	74	)	,
(	74	)	,
(	74	)	,
(	74	)	,
(	74	)	,
(	73	)	,
(	73	)	,
(	73	)	,
(	73	)	,
(	73	)	,
(	73	)	,
(	73	)	,
(	72	)	,
(	72	)	,
(	72	)	,
(	72	)	,
(	72	)	,
(	72	)	,
(	72	)	,
(	71	)	,
(	71	)	,
(	71	)	,
(	71	)	,
(	71	)	,
(	71	)	,
(	71	)	,
(	71	)	,
(	70	)	,
(	70	)	,
(	70	)	,
(	70	)	,
(	70	)	,
(	70	)	,
(	70	)	,
(	69	)	,
(	69	)	,
(	69	)	,
(	69	)	,
(	69	)	,
(	69	)	,
(	69	)	,
(	69	)	,
(	68	)	,
(	68	)	,
(	68	)	,
(	68	)	,
(	68	)	,
(	68	)	,
(	68	)	,
(	68	)	,
(	67	)	,
(	67	)	,
(	67	)	,
(	67	)	,
(	67	)	,
(	67	)	,
(	67	)	,
(	67	)	,
(	66	)	,
(	66	)	,
(	66	)	,
(	66	)	,
(	66	)	,
(	66	)	,
(	66	)	,
(	66	)	,
(	65	)	,
(	65	)	,
(	65	)	,
(	65	)	,
(	65	)	,
(	65	)	,
(	65	)	,
(	65	)	,
(	64	)	,
(	64	)	,
(	64	)	,
(	64	)	,
(	64	)	,
(	64	)	,
(	64	)	,
(	64	)	,
(	64	)	,
(	64	)	,
(	63	)	,
(	63	)	,
(	63	)	,
(	63	)	,
(	63	)	,
(	63	)	,
(	63	)	,
(	63	)	,
(	63	)	,
(	62	)	,
(	62	)	,
(	62	)	,
(	62	)	,
(	62	)	,
(	62	)	,
(	62	)	,
(	62	)	,
(	62	)	,
(	61	)	,
(	61	)	,
(	61	)	,
(	61	)	,
(	61	)	,
(	61	)	,
(	61	)	,
(	61	)	,
(	61	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	10	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	11	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	12	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	13	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	14	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	15	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	16	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	17	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	18	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	19	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	20	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	21	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	22	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	23	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	24	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	25	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	26	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	27	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	28	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	29	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	30	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	31	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	32	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	33	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	34	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	35	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	36	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	37	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	38	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	39	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	40	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	41	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	42	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	43	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	44	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	45	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	46	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	47	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	48	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	49	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	50	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	51	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	52	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	53	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	54	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	55	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	56	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	57	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	58	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	59	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	60	)	,
(	61	)	,
(	61	)	,
(	61	)	,
(	61	)	,
(	62	)	,
(	62	)	,
(	62	)	,
(	62	)	,
(	63	)	,
(	63	)	,
(	63	)	,
(	63	)	,
(	64	)	,
(	64	)	,
(	64	)	,
(	65	)	,
(	65	)	,
(	65	)	,
(	65	)	,
(	66	)	,
(	66	)	,
(	66	)	,
(	66	)	,
(	67	)	,
(	67	)	,
(	67	)	,
(	68	)	,
(	68	)	,
(	68	)	,
(	68	)	,
(	69	)	,
(	69	)	,
(	69	)	,
(	70	)	,
(	70	)	,
(	70	)	,
(	70	)	,
(	71	)	,
(	71	)	,
(	71	)	,
(	72	)	,
(	72	)	,
(	72	)	,
(	72	)	,
(	73	)	,
(	73	)	,
(	73	)	,
(	74	)	,
(	74	)	,
(	74	)	,
(	75	)	,
(	75	)	,
(	75	)	,
(	75	)	,
(	76	)	,
(	76	)	,
(	76	)	,
(	77	)	,
(	77	)	,
(	77	)	,
(	78	)	,
(	78	)	,
(	78	)	,
(	79	)	,
(	79	)	,
(	79	)	,
(	80	)	,
(	80	)	,
(	80	)	,
(	80	)	,
(	81	)	,
(	81	)	,
(	81	)	,
(	82	)	,
(	82	)	,
(	82	)	,
(	83	)	,
(	83	)	,
(	83	)	,
(	84	)	,
(	84	)	,
(	84	)	,
(	85	)	,
(	85	)	,
(	85	)	,
(	86	)	,
(	86	)	,
(	86	)	,
(	87	)	,
(	87	)	,
(	87	)	,
(	88	)	,
(	88	)	,
(	88	)	,
(	89	)	,
(	89	)	,
(	90	)	,
(	90	)	,
(	90	)	,
(	91	)	,
(	91	)	,
(	91	)	,
(	92	)	,
(	92	)	,
(	92	)	,
(	93	)	,
(	93	)	,
(	93	)	,
(	94	)	,
(	94	)	,
(	95	)	,
(	95	)	,
(	95	)	,
(	96	)	,
(	96	)	,
(	96	)	,
(	97	)	,
(	97	)	,
(	97	)	,
(	98	)	,
(	98	)	,
(	99	)	,
(	99	)	,
(	99	)	,
(	100	)	,
(	100	)	,
(	100	)	,
(	101	)	,
(	101	)	,
(	102	)	,
(	102	)	,
(	102	)	,
(	103	)	,
(	103	)	,
(	104	)	,
(	104	)	,
(	104	)	,
(	105	)	,
(	105	)	,
(	105	)	,
(	106	)	,
(	106	)	,
(	107	)	,
(	107	)	,
(	107	)	,
(	108	)	,
(	108	)	,
(	109	)	,
(	109	)	,
(	109	)	,
(	110	)	,
(	110	)	,
(	111	)	,
(	111	)	,
(	112	)	,
(	112	)	,
(	112	)	,
(	113	)	,
(	113	)	,
(	114	)	,
(	114	)	,
(	114	)	,
(	115	)	,
(	115	)	,
(	116	)	,
(	116	)	,
(	117	)	,
(	117	)	,
(	117	)	,
(	118	)	,
(	118	)	,
(	119	)	,
(	119	)	,
(	120	)	,
(	120	)	,
(	120	)	,
(	121	)	,
(	121	)	,
(	122	)	,
(	122	)	,
(	123	)	,
(	123	)	,
(	123	)	,
(	124	)	,
(	124	)	,
(	125	)	,
(	125	)	,
(	126	)	,
(	126	)	,
(	127	)	,
(	127	)	,
(	128	)	,
(	128	)	,
(	128	)	,
(	129	)	,
(	129	)	,
(	130	)	,
(	130	)	,
(	131	)	,
(	131	)	,
(	132	)	,
(	132	)	,
(	133	)	,
(	133	)	,
(	134	)	,
(	134	)	,
(	135	)	,
(	135	)	,
(	135	)	,
(	136	)	,
(	136	)	,
(	137	)	,
(	137	)	,
(	138	)	,
(	138	)	,
(	139	)	,
(	139	)	,
(	140	)	,
(	140	)	,
(	141	)	,
(	141	)	,
(	142	)	,
(	142	)	,
(	143	)	,
(	143	)	,
(	144	)	,
(	144	)	,
(	145	)	,
(	145	)	,
(	146	)	,
(	146	)	,
(	147	)	,
(	147	)	,
(	148	)	,
(	148	)	,
(	149	)	,
(	149	)	,
(	150	)	,
(	150	)	,
(	151	)	,
(	151	)	,
(	152	)	,
(	152	)	,
(	153	)	,
(	153	)	,
(	154	)	,
(	154	)	,
(	155	)	,
(	156	)	,
(	156	)	,
(	157	)	,
(	157	)	,
(	158	)	,
(	158	)	,
(	159	)	,
(	159	)	,
(	160	)	,
(	160	)	,
(	161	)	,
(	161	)	,
(	162	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)	,
(	163	)

);

end package SEVEN_SEG_PWM_LUT;