library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

(8568),
(8548),
(8528),
(8508),
(8488),
(8469),
(8449),
(8430),
(8410),
(8391),
(8371),
(8352),
(8332),
(8313),
(8294),
(8274),
(8255),
(8236),
(8217),
(8198),
(8179),
(8160),
(8141),
(8122),
(8103),
(8084),
(8065),
(8046),
(8027),
(8009),
(7990),
(7971),
(7953),
(7934),
(7916),
(7897),
(7879),
(7860),
(7842),
(7824),
(7805),
(7787),
(7769),
(7751),
(7732),
(7714),
(7696),
(7678),
(7660),
(7642),
(7624),
(7606),
(7588),
(7571),
(7553),
(7535),
(7517),
(7500),
(7482),
(7465),
(7447),
(7429),
(7412),
(7395),
(7377),
(7360),
(7342),
(7325),
(7308),
(7291),
(7273),
(7256),
(7239),
(7222),
(7205),
(7188),
(7171),
(7154),
(7137),
(7120),
(7103),
(7087),
(7070),
(7053),
(7036),
(7020),
(7003),
(6987),
(6970),
(6954),
(6937),
(6921),
(6904),
(6888),
(6872),
(6855),
(6839),
(6823),
(6807),
(6790),
(6774),
(6758),
(6742),
(6726),
(6710),
(6694),
(6678),
(6662),
(6646),
(6631),
(6615),
(6599),
(6583),
(6568),
(6552),
(6536),
(6521),
(6505),
(6490),
(6474),
(6459),
(6443),
(6428),
(6413),
(6397),
(6382),
(6367),
(6352),
(6337),
(6321),
(6306),
(6291),
(6276),
(6261),
(6246),
(6231),
(6216),
(6201),
(6187),
(6172),
(6157),
(6142),
(6128),
(6113),
(6098),
(6084),
(6069),
(6054),
(6040),
(6025),
(6011),
(5997),
(5982),
(5968),
(5953),
(5939),
(5925),
(5911),
(5896),
(5882),
(5868),
(5854),
(5840),
(5826),
(5812),
(5798),
(5784),
(5770),
(5756),
(5742),
(5729),
(5715),
(5701),
(5687),
(5674),
(5660),
(5646),
(5633),
(5619),
(5606),
(5592),
(5579),
(5565),
(5552),
(5538),
(5525),
(5512),
(5498),
(5485),
(5472),
(5459),
(5445),
(5432),
(5419),
(5406),
(5393),
(5380),
(5367),
(5354),
(5341),
(5328),
(5315),
(5303),
(5290),
(5277),
(5264),
(5251),
(5239),
(5226),
(5213),
(5201),
(5188),
(5176),
(5163),
(5151),
(5138),
(5126),
(5113),
(5101),
(5089),
(5076),
(5064),
(5052),
(5040),
(5027),
(5015),
(5003),
(4991),
(4979),
(4967),
(4955),
(4943),
(4931),
(4919),
(4907),
(4895),
(4883),
(4871),
(4859),
(4848),
(4836),
(4824),
(4813),
(4801),
(4789),
(4778),
(4766),
(4754),
(4743),
(4731),
(4720),
(4709),
(4697),
(4686),
(4674),
(4663),
(4652),
(4640),
(4629),
(4618),
(4607),
(4596),
(4584),
(4573),
(4562),
(4551),
(4540),
(4529),
(4518),
(4507),
(4496),
(4485),
(4474),
(4464),
(4453),
(4442),
(4431),
(4420),
(4410),
(4399),
(4388),
(4378),
(4367),
(4356),
(4346),
(4335),
(4325),
(4314),
(4304),
(4293),
(4283),
(4273),
(4262),
(4252),
(4242),
(4231),
(4221),
(4211),
(4201),
(4191),
(4180),
(4170),
(4160),
(4150),
(4140),
(4130),
(4120),
(4110),
(4100),
(4090),
(4080),
(4070),
(4060),
(4051),
(4041),
(4031),
(4021),
(4012),
(4002),
(3992),
(3983),
(3973),
(3963),
(3954),
(3944),
(3935),
(3925),
(3916),
(3906),
(3897),
(3887),
(3878),
(3869),
(3859),
(3850),
(3841),
(3831),
(3822),
(3813),
(3804),
(3794),
(3785),
(3776),
(3767),
(3758),
(3749),
(3740),
(3731),
(3722),
(3713),
(3704),
(3695),
(3686),
(3677),
(3668),
(3660),
(3651),
(3642),
(3633),
(3624),
(3616),
(3607),
(3598),
(3590),
(3581),
(3572),
(3564),
(3555),
(3547),
(3538),
(3530),
(3521),
(3513),
(3504),
(3496),
(3488),
(3479),
(3471),
(3463),
(3454),
(3446),
(3438),
(3430),
(3421),
(3413),
(3405),
(3397),
(3389),
(3381),
(3373),
(3365),
(3357),
(3348),
(3341),
(3333),
(3325),
(3317),
(3309),
(3301),
(3293),
(3285),
(3277),
(3270),
(3262),
(3254),
(3246),
(3239),
(3231),
(3223),
(3216),
(3208),
(3200),
(3193),
(3185),
(3178),
(3170),
(3163),
(3155),
(3148),
(3140),
(3133),
(3125),
(3118),
(3111),
(3103),
(3096),
(3089),
(3081),
(3074),
(3067),
(3060),
(3052),
(3045),
(3038),
(3031),
(3024),
(3017),
(3009),
(3002),
(2995),
(2988),
(2981),
(2974),
(2967),
(2960),
(2953),
(2947),
(2940),
(2933),
(2926),
(2919),
(2912),
(2905),
(2899),
(2892),
(2885),
(2878),
(2872),
(2865),
(2858),
(2852),
(2845),
(2839),
(2832),
(2825),
(2819),
(2812),
(2806),
(2799),
(2793),
(2786),
(2780),
(2773),
(2767),
(2761),
(2754),
(2748),
(2742),
(2735),
(2729),
(2723),
(2716),
(2710),
(2704),
(2698),
(2692),
(2685),
(2679),
(2673),
(2667),
(2661),
(2655),
(2649),
(2643),
(2637),
(2631),
(2625),
(2619),
(2613),
(2607),
(2601),
(2595),
(2589),
(2583),
(2577),
(2571),
(2566),
(2560),
(2554),
(2548),
(2542),
(2537),
(2531),
(2525),
(2520),
(2514),
(2508),
(2503),
(2497),
(2491),
(2486),
(2480),
(2475),
(2469),
(2464),
(2458),
(2453),
(2447),
(2442),
(2436),
(2431),
(2425),
(2420),
(2415),
(2409),
(2404),
(2398),
(2393),
(2388),
(2383),
(2377),
(2372),
(2367),
(2362),
(2356),
(2351),
(2346),
(2341),
(2336),
(2331),
(2325),
(2320),
(2315),
(2310),
(2305),
(2300),
(2295),
(2290),
(2285),
(2280),
(2275),
(2270),
(2265),
(2260),
(2256),
(2251),
(2246),
(2241),
(2236),
(2231),
(2226),
(2222),
(2217),
(2212),
(2207),
(2203),
(2198),
(2193),
(2189),
(2184),
(2179),
(2175),
(2170),
(2165),
(2161),
(2156),
(2151),
(2147),
(2142),
(2138),
(2133),
(2129),
(2124),
(2120),
(2115),
(2111),
(2107),
(2102),
(2098),
(2093),
(2089),
(2085),
(2080),
(2076),
(2072),
(2067),
(2063),
(2059),
(2054),
(2050),
(2046),
(2042),
(2037),
(2033),
(2029),
(2025),
(2021),
(2017),
(2012),
(2008),
(2004),
(2000),
(1996),
(1992),
(1988),
(1984),
(1980),
(1976),
(1972),
(1968),
(1964),
(1960),
(1956),
(1952),
(1948),
(1944),
(1940),
(1936),
(1932),
(1928),
(1925),
(1921),
(1917),
(1913),
(1909),
(1906),
(1902),
(1898),
(1894),
(1890),
(1887),
(1883),
(1879),
(1876),
(1872),
(1868),
(1865),
(1861),
(1857),
(1854),
(1850),
(1847),
(1843),
(1839),
(1836),
(1832),
(1829),
(1825),
(1822),
(1818),
(1815),
(1811),
(1808),
(1804),
(1801),
(1797),
(1794),
(1791),
(1787),
(1784),
(1780),
(1777),
(1774),
(1770),
(1767),
(1764),
(1760),
(1757),
(1754),
(1750),
(1747),
(1744),
(1741),
(1737),
(1734),
(1731),
(1728),
(1725),
(1721),
(1718),
(1715),
(1712),
(1709),
(1706),
(1703),
(1699),
(1696),
(1693),
(1690),
(1687),
(1684),
(1681),
(1678),
(1675),
(1672),
(1669),
(1666),
(1663),
(1660),
(1657),
(1654),
(1651),
(1648),
(1645),
(1642),
(1639),
(1637),
(1634),
(1631),
(1628),
(1625),
(1622),
(1619),
(1617),
(1614),
(1611),
(1608),
(1605),
(1603),
(1600),
(1597),
(1594),
(1592),
(1589),
(1586),
(1584),
(1581),
(1578),
(1575),
(1573),
(1570),
(1567),
(1565),
(1562),
(1560),
(1557),
(1554),
(1552),
(1549),
(1547),
(1544),
(1541),
(1539),
(1536),
(1534),
(1531),
(1529),
(1526),
(1524),
(1521),
(1519),
(1516),
(1514),
(1511),
(1509),
(1507),
(1504),
(1502),
(1499),
(1497),
(1494),
(1492),
(1490),
(1487),
(1485),
(1483),
(1480),
(1478),
(1476),
(1473),
(1471),
(1469),
(1466),
(1464),
(1462),
(1460),
(1457),
(1455),
(1453),
(1451),
(1448),
(1446),
(1444),
(1442),
(1440),
(1437),
(1435),
(1433),
(1431),
(1429),
(1427),
(1424),
(1422),
(1420),
(1418),
(1416),
(1414),
(1412),
(1410),
(1407),
(1405),
(1403),
(1401),
(1399),
(1397),
(1395),
(1393),
(1391),
(1389),
(1387),
(1385),
(1383),
(1381),
(1379),
(1377),
(1375),
(1373),
(1371),
(1369),
(1367),
(1365),
(1364),
(1362),
(1360),
(1358),
(1356),
(1354),
(1352),
(1350),
(1348),
(1347),
(1345),
(1343),
(1341),
(1339),
(1337),
(1335),
(1334),
(1332),
(1330),
(1328),
(1326),
(1325),
(1323),
(1321),
(1319),
(1318),
(1316),
(1314),
(1312),
(1311),
(1309),
(1307),
(1305),
(1304),
(1302),
(1300),
(1299),
(1297),
(1295),
(1294),
(1292),
(1290),
(1289),
(1287),
(1285),
(1284),
(1282),
(1281),
(1279),
(1277),
(1276),
(1274),
(1272),
(1271),
(1269),
(1268),
(1266),
(1265),
(1263),
(1261),
(1260),
(1258),
(1257),
(1255),
(1254),
(1252),
(1251),
(1249),
(1248),
(1246),
(1245),
(1243),
(1242),
(1240),
(1239),
(1237),
(1236),
(1234),
(1233),
(1232),
(1230),
(1229),
(1227),
(1226),
(1224),
(1223),
(1222),
(1220),
(1219),
(1217),
(1216),
(1215),
(1213),
(1212),
(1210),
(1209),
(1208),
(1206),
(1205),
(1204),
(1202),
(1201),
(1200),
(1198),
(1197),
(1196),
(1194),
(1193),
(1192),
(1190),
(1189),
(1188),
(1187),
(1185),
(1184),
(1183),
(1181),
(1180),
(1179),
(1178),
(1176),
(1175),
(1174),
(1173),
(1171),
(1170),
(1169),
(1168),
(1167),
(1165),
(1164),
(1163),
(1162),
(1161),
(1159),
(1158),
(1157),
(1156),
(1155),
(1153),
(1152),
(1151),
(1150),
(1149),
(1148),
(1146),
(1145),
(1144),
(1143),
(1142),
(1141),
(1140),
(1139),
(1137),
(1136),
(1135),
(1134),
(1133),
(1132),
(1131),
(1130),
(1129),
(1128),
(1126),
(1125),
(1124),
(1123),
(1122),
(1121),
(1120),
(1119),
(1118),
(1117),
(1116),
(1115),
(1114),
(1113),
(1112),
(1111),
(1110),
(1109),
(1108),
(1107),
(1106),
(1104),
(1103),
(1102),
(1101),
(1100),
(1099),
(1098),
(1097),
(1097),
(1096),
(1095),
(1094),
(1093),
(1092),
(1091),
(1090),
(1089),
(1088),
(1087),
(1086),
(1085),
(1084),
(1083),
(1082),
(1081),
(1080),
(1079),
(1078),
(1077),
(1076),
(1075),
(1075),
(1074),
(1073),
(1072),
(1071),
(1070),
(1069),
(1068),
(1067),
(1066),
(1065),
(1065),
(1064),
(1063),
(1062),
(1061),
(1060),
(1059),
(1058),
(1058),
(1057),
(1056),
(1055),
(1054),
(1053),
(1052),
(1051),
(1051),
(1050),
(1049),
(1048),
(1047),
(1046),
(1045),
(1045),
(1044),
(1043),
(1042),
(1041),
(1040),
(1040),
(1039),
(1038),
(1037),
(1036),
(1036),
(1035),
(1034),
(1033),
(1032),
(1031),
(1031),
(1030),
(1029),
(1028),
(1027),
(1027),
(1026),
(1025),
(1024),
(1023),
(1023),
(1022),
(1021),
(1020),
(1020),
(1019),
(1018),
(1017),
(1016),
(1016),
(1015),
(1014),
(1013),
(1013),
(1012),
(1011),
(1010),
(1009),
(1009),
(1008),
(1007),
(1006),
(1006),
(1005),
(1004),
(1003),
(1003),
(1002),
(1001),
(1000),
(1000),
(999),
(998),
(997),
(997),
(996),
(995),
(995),
(994),
(993),
(992),
(992),
(991),
(990),
(989),
(989),
(988),
(987),
(986),
(986),
(985),
(984),
(984),
(983),
(982),
(981),
(981),
(980),
(979),
(979),
(978),
(977),
(976),
(976),
(975),
(974),
(974),
(973),
(972),
(972),
(971),
(970),
(969),
(969),
(968),
(967),
(967),
(966),
(965),
(965),
(964),
(963),
(962),
(962),
(961),
(960),
(960),
(959),
(958),
(958),
(957),
(956),
(956),
(955),
(954),
(954),
(953),
(952),
(951),
(951),
(950),
(949),
(949),
(948),
(947),
(947),
(946),
(945),
(945),
(944),
(943),
(943),
(942),
(941),
(941),
(940),
(939),
(939),
(938),
(937),
(937),
(936),
(935),
(935),
(934),
(933),
(933),
(932),
(931),
(931),
(930),
(929),
(929),
(928),
(927),
(927),
(926),
(925),
(924),
(924),
(923),
(922),
(922),
(921),
(920),
(920),
(919),
(918),
(918),
(917),
(916),
(916),
(915),
(914),
(914),
(913),
(912),
(912),
(911),
(910),
(910),
(909),
(908),
(908),
(907),
(906),
(906),
(905),
(904),
(904),
(903),
(902),
(902),
(901),
(900),
(900),
(899),
(898),
(898),
(897),
(896),
(896),
(895),
(894),
(894),
(893),
(892),
(892),
(891),
(890),
(890),
(889),
(888),
(888),
(887),
(886),
(886),
(885),
(884),
(884),
(883),
(882),
(882),
(881),
(880),
(880),
(879),
(878),
(878),
(877),
(876),
(876),
(875),
(874),
(873),
(873),
(872),
(871),
(871),
(870),
(869),
(869),
(868),
(867),
(867),
(866),
(865),
(865),
(864),
(863),
(863),
(862),
(861),
(860),
(860),
(859),
(858),
(858),
(857),
(856),
(856),
(855),
(854),
(854),
(853),
(852),
(851),
(851),
(850),
(849),
(849),
(848),
(847),
(847),
(846),
(845),
(844),
(844),
(843),
(842),
(842),
(841),
(840),
(839),
(839),
(838),
(837),
(837),
(836),
(835),
(835),
(834),
(833),
(832),
(832),
(831),
(830),
(829),
(829),
(828),
(827),
(827),
(826),
(825),
(824),
(824),
(823),
(822),
(822),
(821),
(820),
(819),
(819),
(818),
(817),
(816),
(816),
(815),
(814),
(814),
(813),
(812),
(811),
(811),
(810),
(809),
(808),
(808),
(807),
(806),
(805),
(805),
(804),
(803),
(802),
(802),
(801),
(800),
(799),
(799),
(798),
(797),
(796),
(796),
(795),
(794),
(793),
(793),
(792),
(791),
(790),
(790),
(789),
(788),
(787),
(787),
(786),
(785),
(784),
(783),
(783),
(782),
(781),
(780),
(780),
(779),
(778),
(777),
(776),
(776),
(775),
(774),
(773),
(773),
(772),
(771),
(770),
(769),
(769),
(768),
(767),
(766),
(765),
(765),
(764),
(763),
(762),
(762),
(761),
(760),
(759),
(758),
(758),
(757),
(756),
(755),
(754),
(754),
(753),
(752),
(751),
(750),
(750),
(749),
(748),
(747),
(746),
(745),
(745),
(744),
(743),
(742),
(741),
(741),
(740),
(739),
(738),
(737),
(736),
(736),
(735),
(734),
(733),
(732),
(731),
(731),
(730),
(729),
(728),
(727),
(726),
(726),
(725),
(724),
(723),
(722),
(721),
(721),
(720),
(719),
(718),
(717),
(716),
(716),
(715),
(714),
(713),
(712),
(711),
(710),
(710),
(709),
(708),
(707),
(706),
(705),
(704),
(704),
(703),
(702),
(701),
(700),
(699),
(698),
(698),
(697),
(696),
(695),
(694),
(693),
(692),
(691),
(691),
(690),
(689),
(688),
(687),
(686),
(685),
(684),
(684),
(683),
(682),
(681),
(680),
(679),
(678),
(677),
(677),
(676),
(675),
(674),
(673),
(672),
(671),
(670),
(669),
(669),
(668),
(667),
(666),
(665),
(664),
(663),
(662),
(661),
(661),
(660),
(659),
(658),
(657),
(656),
(655),
(654),
(653),
(652),
(651),
(651),
(650),
(649),
(648),
(647),
(646),
(645),
(644),
(643),
(642),
(641),
(641),
(640),
(639),
(638),
(637),
(636),
(635),
(634),
(633),
(632),
(631),
(630),
(630),
(629),
(628),
(627),
(626),
(625),
(624),
(623),
(622),
(621),
(620),
(619),
(618),
(618),
(617),
(616),
(615),
(614),
(613),
(612),
(611),
(610),
(609),
(608),
(607),
(606),
(605),
(604),
(604),
(603),
(602),
(601),
(600),
(599),
(598),
(597),
(596),
(595),
(594),
(593),
(592),
(591),
(590),
(589),
(589),
(588),
(587),
(586),
(585),
(584),
(583),
(582),
(581),
(580),
(579),
(578),
(577),
(576),
(575),
(574),
(573),
(572),
(572),
(571),
(570),
(569),
(568),
(567),
(566),
(565),
(564),
(563),
(562),
(561),
(560),
(559),
(558),
(557),
(556),
(555),
(554),
(554),
(553),
(552),
(551),
(550),
(549),
(548),
(547),
(546),
(545),
(544),
(543),
(542),
(541),
(540),
(539),
(538),
(537),
(536),
(535),
(535),
(534),
(533),
(532),
(531),
(530),
(529),
(528),
(527),
(526),
(525),
(524),
(523),
(522),
(521),
(520),
(519),
(518),
(518),
(517),
(516),
(515),
(514),
(513),
(512),
(511),
(510),
(509),
(508),
(507),
(506),
(505),
(504),
(503),
(502),
(501),
(501),
(500),
(499),
(498),
(497),
(496),
(495),
(494),
(493),
(492),
(491),
(490),
(489),
(488),
(487),
(487),
(486),
(485),
(484),
(483),
(482),
(481),
(480),
(479),
(478),
(477),
(476),
(475),
(475),
(474),
(473),
(472),
(471),
(470),
(469),
(468),
(467),
(466),
(465),
(464),
(464),
(463),
(462),
(461),
(460),
(459),
(458),
(457),
(456),
(455),
(454),
(454),
(453),
(452),
(451),
(450),
(449),
(448),
(447),
(446),
(445),
(445),
(444),
(443),
(442),
(441),
(440),
(439),
(438),
(438),
(437),
(436),
(435),
(434),
(433),
(432),
(431),
(431),
(430),
(429),
(428),
(427),
(426),
(425),
(424),
(424),
(423),
(422),
(421),
(420),
(419),
(418),
(418),
(417),
(416),
(415),
(414),
(413),
(413),
(412),
(411),
(410),
(409),
(408),
(408),
(407),
(406),
(405),
(404),
(403),
(403),
(402),
(401),
(400),
(399),
(399),
(398),
(397),
(396),
(395),
(394),
(394),
(393),
(392),
(391),
(391),
(390),
(389),
(388),
(387),
(387),
(386),
(385),
(384),
(383),
(383),
(382),
(381),
(380),
(380),
(379),
(378),
(377),
(377),
(376),
(375),
(374),
(374),
(373),
(372),
(371),
(371),
(370),
(369),
(368),
(368),
(367),
(366),
(366),
(365),
(364),
(363),
(363),
(362),
(361),
(361),
(360),
(359),
(359),
(358),
(357),
(356),
(356),
(355),
(354),
(354),
(353),
(352),
(352),
(351),
(350),
(350),
(349),
(349),
(348),
(347),
(347),
(346),
(345),
(345),
(344),
(343),
(343),
(342),
(342),
(341),
(340),
(340),
(339),
(339),
(338),
(337),
(337),
(336),
(336),
(335),
(334),
(334),
(333),
(333),
(332),
(332),
(331),
(330),
(330),
(329),
(329),
(328),
(328),
(327),
(327),
(326),
(326),
(325),
(325),
(324),
(324),
(323),
(322),
(322),
(321),
(321),
(321),
(320),
(320),
(319),
(319),
(318),
(318),
(317),
(317),
(316),
(316),
(315),
(315),
(315),
(314),
(314),
(313),
(313),
(312),
(312),
(312),
(311),
(311),
(310),
(310),
(310),
(309),
(309),
(308),
(308),
(308),
(307),
(307),
(307),
(306),
(306),
(306),
(305),
(305),
(305),
(304),
(304),
(304),
(303),
(303),
(303),
(302),
(302),
(302),
(302),
(301),
(301),
(301),
(301),
(300),
(300),
(300),
(300),
(299),
(299),
(299),
(299),
(298),
(298),
(298),
(298),
(298),
(297),
(297),
(297),
(297),
(297),
(296),
(296),
(296),
(296),
(296),
(296),
(296),
(295),
(295),
(295),
(295),
(295),
(295),
(295),
(295),
(295),
(295),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(294),
(295),
(295),
(295),
(295),
(295),
(295),
(295),
(295),
(295),
(296),
(296),
(296),
(296),
(296),
(296),
(297),
(297),
(297),
(297),
(297),
(298),
(298),
(298),
(298),
(298),
(299),
(299),
(299),
(299),
(300),
(300),
(300),
(301),
(301),
(301),
(301),
(302),
(302),
(302),
(303),
(303),
(303),
(304),
(304),
(305),
(305),
(305),
(306),
(306),
(307),
(307),
(307),
(308),
(308),
(309),
(309),
(310),
(310),
(311),
(311),
(312),
(312),
(313),
(313),
(314),
(314),
(315),
(315),
(316),
(316),
(317),
(318),
(318),
(319),
(319),
(320),
(321),
(321),
(322),
(322),
(323),
(324),
(324),
(325),
(326),
(326),
(327),
(328),
(329),
(329),
(330),
(331),
(331),
(332),
(333),
(334),
(335),
(335),
(336),
(337),
(338),
(339),
(339),
(340),
(341),
(342),
(343),
(344),
(345),
(346),
(346),
(347),
(348),
(349),
(350),
(351),
(352),
(353),
(354),
(355),
(356),
(357),
(358),
(359),
(360),
(361),
(362),
(363),
(364),
(365),
(366),
(367),
(369),
(370),
(371),
(372),
(373),
(374),
(375),
(377),
(378),
(379),
(380),
(381),
(383),
(384),
(385),
(386),
(388),
(389),
(390),
(391),
(393),
(394),
(395),
(397),
(398),
(399),
(401),
(402),
(403),
(405),
(406),
(408),
(409),
(411),
(412),
(413),
(415),
(416),
(418),
(419),
(421),
(422),
(424),
(425),
(427),
(429),
(430),
(432),
(433),
(435),
(437),
(438),
(440),
(441),
(443),
(445),
(446),
(448),
(450),
(452),
(453),
(455),
(457),
(459),
(460),
(462),
(464),
(466),
(467),
(469),
(471),
(473),
(475),
(477),
(479),
(480),
(482),
(484),
(486),
(488),
(490),
(492),
(494),
(496),
(498),
(500),
(502),
(504),
(506),
(508),
(510),
(512),
(515),
(517),
(519),
(521),
(523),
(525),
(527),
(530),
(532),
(534),
(536),
(538),
(541),
(543),
(545),
(547),
(550),
(552),
(554),
(557),
(559),
(561),
(564),
(566),
(569),
(571),
(573),
(576),
(578),
(581),
(583),
(586),
(588),
(591),
(593),
(596),
(598),
(601),
(604),
(606),
(609),
(611),
(614),
(617),
(619),
(622),
(625),
(627),
(630),
(633),
(636),
(638),
(641),
(644),
(647),
(649),
(652),
(655),
(658),
(661),
(664),
(667),
(670),
(672),
(675),
(678),
(681),
(684),
(687),
(690),
(693),
(696),
(699),
(703),
(706),
(709),
(712),
(715),
(718),
(721),
(724),
(728),
(731),
(734),
(737),
(740),
(744),
(747),
(750),
(754),
(757),
(760),
(764),
(767),
(770),
(774),
(777),
(781),
(784),
(787),
(791),
(794),
(798),
(801),
(805),
(809),
(812),
(816),
(819),
(823),
(827),
(830),
(834),
(838),
(841),
(845),
(849),
(852),
(856),
(860),
(864),
(868),
(871),
(875),
(879),
(883),
(887),
(891),
(895),
(899),
(902),
(906),
(910),
(914),
(918),
(922),
(927),
(931),
(935),
(939),
(943),
(947),
(951),
(955),
(960),
(964),
(968),
(972),
(976),
(981),
(985),
(989),
(994),
(998),
(1002),
(1007),
(1011),
(1016),
(1020),
(1024),
(1029),
(1033),
(1038),
(1042),
(1047),
(1051),
(1056),
(1061),
(1065),
(1070),
(1074),
(1079),
(1084),
(1088),
(1093),
(1098),
(1103),
(1107),
(1112),
(1117),
(1122),
(1127),
(1132),
(1136),
(1141),
(1146),
(1151),
(1156),
(1161),
(1166),
(1171),
(1176),
(1181),
(1186),
(1191),
(1196),
(1201),
(1207),
(1212),
(1217),
(1222),
(1227),
(1233),
(1238),
(1243),
(1248),
(1254),
(1259),
(1264),
(1270),
(1275),
(1281),
(1286),
(1291),
(1297),
(1302),
(1308),
(1313),
(1319),
(1324),
(1330),
(1336),
(1341),
(1347),
(1353),
(1358),
(1364),
(1370),
(1375),
(1381),
(1387),
(1393),
(1399),
(1404),
(1410),
(1416),
(1422),
(1428),
(1434),
(1440),
(1446),
(1452),
(1458),
(1464),
(1470),
(1476),
(1482),
(1488),
(1495),
(1501),
(1507),
(1513),
(1519),
(1526),
(1532),
(1538),
(1545),
(1551),
(1557),
(1564),
(1570),
(1576),
(1583),
(1589),
(1596),
(1602),
(1609),
(1615),
(1622),
(1629),
(1635),
(1642),
(1649),
(1655),
(1662),
(1669),
(1675),
(1682),
(1689),
(1696),
(1703),
(1710),
(1716),
(1723),
(1730),
(1737),
(1744),
(1751),
(1758),
(1765),
(1772),
(1779),
(1787),
(1794),
(1801),
(1808),
(1815),
(1823),
(1830),
(1837),
(1844),
(1852),
(1859),
(1866),
(1874),
(1881),
(1889),
(1896),
(1904),
(1911),
(1919),
(1926),
(1934),
(1941),
(1949),
(1957),
(1964),
(1972),
(1980),
(1987),
(1995),
(2003),
(2011),
(2019),
(2026),
(2034),
(2042),
(2050),
(2058),
(2066),
(2074),
(2082),
(2090),
(2098),
(2106),
(2115),
(2123),
(2131),
(2139),
(2147),
(2156),
(2164),
(2172),
(2180),
(2189),
(2197),
(2206),
(2214),
(2222),
(2231),
(2239),
(2248),
(2257),
(2265),
(2274),
(2282),
(2291),
(2300),
(2308),
(2317),
(2326),
(2335),
(2343),
(2352),
(2361),
(2370),
(2379),
(2388),
(2397),
(2406),
(2415),
(2424),
(2433),
(2442),
(2451),
(2460),
(2469),
(2479),
(2488),
(2497),
(2506),
(2516),
(2525),
(2534),
(2544),
(2553),
(2563),
(2572),
(2582),
(2591),
(2601),
(2610),
(2620),
(2629),
(2639),
(2649),
(2659),
(2668),
(2678),
(2688),
(2698),
(2707),
(2717),
(2727),
(2737),
(2747),
(2757),
(2767),
(2777),
(2787),
(2797),
(2807),
(2818),
(2828),
(2838),
(2848),
(2858),
(2869),
(2879),
(2889),
(2900),
(2910),
(2921),
(2931),
(2942),
(2952),
(2963),
(2973),
(2984),
(2994),
(3005),
(3016),
(3027),
(3037),
(3048),
(3059),
(3070),
(3081),
(3091),
(3102),
(3113),
(3124),
(3135),
(3146),
(3157),
(3168),
(3180),
(3191),
(3202),
(3213),
(3224),
(3236),
(3247),
(3258),
(3270),
(3281),
(3293),
(3304),
(3315),
(3327),
(3339),
(3350),
(3362),
(3373),
(3385),
(3397),
(3408),
(3420),
(3432),
(3444),
(3456),
(3468),
(3479),
(3491),
(3503),
(3515),
(3527),
(3539),
(3552),
(3564),
(3576),
(3588),
(3600),
(3612),
(3625),
(3637),
(3649),
(3662),
(3674),
(3687),
(3699),
(3712),
(3724),
(3737),
(3749),
(3762),
(3775),
(3787),
(3800),
(3813),
(3826),
(3838),
(3851),
(3864),
(3877),
(3890),
(3903),
(3916),
(3929),
(3942),
(3955),
(3968),
(3982),
(3995),
(4008),
(4021),
(4035),
(4048),
(4061),
(4075),
(4088),
(4102),
(4115),
(4129),
(4142),
(4156),
(4170),
(4183),
(4197),
(4211),
(4225),
(4238),
(4252),
(4266),
(4280),
(4294),
(4308),
(4322),
(4336),
(4350),
(4364),
(4378),
(4393),
(4407),
(4421),
(4435),
(4450),
(4464),
(4478),
(4493),
(4507),
(4522),
(4536),
(4551),
(4566),
(4580),
(4595),
(4610),
(4624),
(4639),
(4654),
(4669),
(4684),
(4698),
(4713),
(4728),
(4743),
(4759),
(4774),
(4789),
(4804),
(4819),
(4834),
(4850),
(4865),
(4880),
(4896),
(4911),
(4927),
(4942),
(4958),
(4973),
(4989),
(5004),
(5020),
(5036),
(5051),
(5067),
(5083),
(5099),
(5115),
(5131),
(5147),
(5163),
(5179),
(5195),
(5211),
(5227),
(5243),
(5259),
(5276),
(5292),
(5308),
(5325),
(5341),
(5358),
(5374),
(5391),
(5407),
(5424),
(5440),
(5457),
(5474),
(5490),
(5507),
(5524),
(5541),
(5558),
(5575),
(5592),
(5609),
(5626),
(5643),
(5660),
(5677),
(5694),
(5712),
(5729),
(5746),
(5764),
(5781),
(5798),
(5816),
(5833),
(5851),
(5869),
(5886),
(5904),
(5922),
(5939),
(5957),
(5975),
(5993),
(6011),
(6029),
(6047),
(6065),
(6083),
(6101),
(6119),
(6137),
(6155),
(6174),
(6192),
(6210),
(6229),
(6247),
(6266),
(6284),
(6303),
(6321),
(6340),
(6359),
(6377),
(6396),
(6415),
(6434),
(6453),
(6472),
(6490),
(6509),
(6529),
(6548),
(6567),
(6586),
(6605),
(6624),
(6644),
(6663),
(6682),
(6702),
(6721),
(6741),
(6760),
(6780),
(6799),
(6819),
(6839),
(6858),
(6878),
(6898),
(6918),
(6938),
(6958),
(6978),
(6998),
(7018),
(7038),
(7058),
(7078),
(7099),
(7119),
(7139),
(7160),
(7180),
(7201),
(7221),
(7242),
(7262),
(7283),
(7304),
(7324),
(7345),
(7366),
(7387),
(7408),
(7429),
(7450),
(7471),
(7492),
(7513),
(7534),
(7555),
(7576),
(7598),
(7619),
(7640),
(7662),
(7683),
(7705),
(7726),
(7748),
(7770),
(7791),
(7813),
(7835),
(7857),
(7879),
(7900),
(7922),
(7944),
(7967),
(7989),
(8011),
(8033),
(8055),
(8077),
(8100),
(8122),
(8145),
(8167),
(8190),
(8212),
(8235),
(8257),
(8280),
(8303),
(8326),
(8348),
(8371),
(8394),
(8417),
(8440),
(8463),
(8486),
(8509),
(8533),
(8556),
(8579),
(8602),
(8626),
(8649),
(8673),
(8696),
(8720),
(8743),
(8767),
(8791),
(8815),
(8838),
(8862),
(8886),
(8910),
(8934),
(8958),
(8982),
(9006),
(9031),
(9055),
(9079),
(9103),
(9128),
(9152),
(9177),
(9201),
(9226),
(9250),
(9275),
(9300),
(9325),
(9349),
(9374),
(9399),
(9424),
(9449),
(9474),
(9499),
(9524),
(9550),
(9575),
(9600),
(9625),
(9651),
(9676),
(9702),
(9727),
(9753),
(9779),
(9804),
(9830),
(9856),
(9882),
(9908),
(9933),
(9959),
(9986),
(10012),
(10038),
(10064),
(10090),
(10116),
(10143),
(10169),
(10196),
(10222),
(10249),
(10275),
(10302),
(10329),
(10355),
(10382),
(10409),
(10436),
(10463),
(10490),
(10517),
(10544),
(10571),
(10598),
(10626),
(10653),
(10680),
(10708),
(10735),
(10763),
(10790),
(10818),
(10846),
(10873),
(10901),
(10929),
(10957),
(10985),
(11013),
(11041),
(11069),
(11097),
(11125),
(11154),
(11182),
(11210),
(11239),
(11267),
(11296),
(11324),
(11353),
(11381),
(11410),
(11439),
(11468),
(11497),
(11526),
(11555),
(11584),
(11613),
(11642),
(11671),
(11700),
(11730),
(11759),
(11788),
(11818),
(11848),
(11877),
(11907),
(11936),
(11966),
(11996),
(12026),
(12056),
(12086),
(12116),
(12146),
(12176),
(12206),
(12236),
(12267),
(12297),
(12327),
(12358),
(12388),
(12419),
(12450),
(12480),
(12511),
(12542),
(12573),
(12604),
(12635),
(12666),
(12697),
(12728),
(12759),
(12790),
(12822),
(12853),
(12884),
(12916),
(12947),
(12979),
(13011),
(13042),
(13074),
(13106),
(13138),
(13170),
(13202),
(13234),
(13266),
(13298),
(13330),
(13362),
(13395),
(13427),
(13459),
(13492),
(13525),
(13557),
(13590),
(13623),
(13655),
(13688),
(13721),
(13754),
(13787),
(13820),
(13853),
(13886),
(13920),
(13953),
(13986),
(14020),
(14053),
(14087),
(14120),
(14154),
(14188),
(14222),
(14255),
(14289),
(14323),
(14357),
(14391),
(14425),
(14460),
(14494),
(14528),
(14563),
(14597),
(14632),
(14666),
(14701),
(14735),
(14770),
(14805),
(14840),
(14875),
(14910),
(14945),
(14980),
(15015),
(15050),
(15085),
(15121),
(15156),
(15192),
(15227),
(15263),
(15298),
(15334),
(15370),
(15406),
(15442),
(15477),
(15514),
(15550),
(15586),
(15622),
(15658),
(15694),
(15731),
(15767),
(15804),
(15840),
(15877),
(15914),
(15950),
(15987),
(16024),
(16061),
(16098),
(16135),
(16172),
(16209),
(16247),
(16284),
(16321),
(16359),
(16396),
(16434),
(16472),
(16509),
(16547),
(16585),
(16623),
(16661),
(16699),
(16737),
(16775),
(16813),
(16851),
(16890),
(16928),
(16967),
(17005),
(17044),
(17082),
(17121),
(17160),
(17199),
(17238),
(17277),
(17316),
(17355),
(17394),
(17433),
(17472),
(17512),
(17551),
(17591),
(17630),
(17670),
(17710),
(17749),
(17789),
(17829),
(17869),
(17909),
(17949),
(17989),
(18030),
(18070),
(18110),
(18151),
(18191),
(18232),
(18272),
(18313),
(18354),
(18394),
(18435),
(18476),
(18517),
(18558),
(18600),
(18641),
(18682),
(18723),
(18765),
(18806),
(18848),
(18890),
(18931),
(18973),
(19015),
(19057),
(19099),
(19141),
(19183),
(19225),
(19267),
(19309),
(19352),
(19394),
(19437),
(19479),
(19522),
(19565),
(19607),
(19650),
(19693),
(19736),
(19779),
(19822),
(19866),
(19909),
(19952),
(19996),
(20039),
(20083),
(20126),
(20170),
(20214),
(20257),
(20301),
(20345),
(20389),
(20433),
(20478),
(20522),
(20566),
(20611),
(20655),
(20700),
(20744),
(20789),
(20834),
(20878),
(20923),
(20968),
(21013),
(21058),
(21103),
(21149),
(21194),
(21239),
(21285),
(21330),
(21376),
(21422),
(21467),
(21513),
(21559),
(21605),
(21651),
(21697),
(21743),
(21789),
(21836),
(21882),
(21929),
(21975),
(22022),
(22068),
(22115),
(22162),
(22209),
(22256),
(22303),
(22350),
(22397),
(22444),
(22492),
(22539),
(22587),
(22634),
(22682),
(22729),
(22777),
(22825),
(22873),
(22921),
(22969),
(23017),
(23065),
(23114),
(23162),
(23210),
(23259),
(23307),
(23356),
(23405),
(23454),
(23503),
(23552),
(23601),
(23650),
(23699),
(23748),
(23797),
(23847),
(23896),
(23946),
(23996),
(24045),
(24095),
(24145),
(24195),
(24245),
(24295),
(24345),
(24395),
(24446),
(24496),
(24547),
(24597),
(24648),
(24698),
(24749),
(24800),
(24851),
(24902),
(24953),
(25004),
(25056),
(25107),
(25158),
(25210),
(25261),
(25313),
(25365),
(25416),
(25468),
(25520),
(25572),
(25624),
(25677),
(25729),
(25781),
(25834),
(25886),
(25939),
(25991),
(26044),
(26097),
(26150),
(26203),
(26256),
(26309),
(26362),
(26415),
(26469),
(26522),
(26576),
(26629),
(26683),
(26737),
(26790),
(26844),
(26898),
(26952),
(27007),
(27061),
(27115),
(27169),
(27224),
(27279),
(27333),
(27388),
(27443),
(27498),
(27553),
(27608),
(27663),
(27718),
(27773),
(27829),
(27884),
(27939),
(27995),
(28051),
(28107),
(28162),
(28218),
(28274),
(28330),
(28387),
(28443),
(28499),
(28556),
(28612),
(28669),
(28725),
(28782),
(28839),
(28896),
(28953),
(29010),
(29067),
(29124),
(29182),
(29239),
(29297),
(29354),
(29412),
(29470),
(29528),
(29585),
(29643),
(29702),
(29760),
(29818),
(29876),
(29935),
(29993),
(30052),
(30111),
(30169),
(30228),
(30287),
(30346),
(30405),
(30464),
(30524),
(30583),
(30642),
(30702),
(30762),
(30821),
(30881),
(30941),
(31001),
(31061),
(31121),
(31181),
(31241),
(31302),
(31362),
(31423),
(31484),
(31544),
(31605),
(31666),
(31727),
(31788),
(31849),
(31910),
(31972),
(32033),
(32095),
(32156),
(32218),
(32280),
(32341),
(32403),
(32465),
(32528),
(32590),
(32652),
(32714),
(32777),
(32839),
(32902),
(32965),
(33028),
(33091),
(33154),
(33217),
(33280),
(33343),
(33406),
(33470),
(33533),
(33597),
(33661),
(33724),
(33788),
(33852),
(33916),
(33981),
(34045),
(34109),
(34173),
(34238),
(34303),
(34367),
(34432),
(34497),
(34562),
(34627),
(34692),
(34757),
(34823),
(34888),
(34953),
(35019),
(35085),
(35151),
(35216),
(35282),
(35348),
(35415),
(35481),
(35547),
(35613),
(35680),
(35747),
(35813),
(35880),
(35947),
(36014),
(36081),
(36148),
(36215),
(36283),
(36350),
(36418),
(36485),
(36553),
(36621),
(36688),
(36756),
(36825),
(36893),
(36961),
(37029),
(37098),
(37166),
(37235),
(37304),
(37372),
(37441),
(37510),
(37579),
(37649),
(37718),
(37787),
(37857),
(37926),
(37996),
(38066),
(38136),
(38205),
(38276),
(38346),
(38416),
(38486),
(38557),
(38627),
(38698),
(38768),
(38839),
(38910),
(38981),
(39052),
(39123),
(39195),
(39266),
(39337),
(39409),
(39481),
(39552),
(39624),
(39696),
(39768),
(39840),
(39913),
(39985),
(40057),
(40130),
(40203),
(40275),
(40348),
(40421),
(40494),
(40567),
(40640),
(40714),
(40787),
(40861),
(40934),
(41008),
(41082),
(41156),
(41230),
(41304),
(41378),
(41452),
(41526),
(41601),
(41676),
(41750),
(41825),
(41900),
(41975),
(42050),
(42125),
(42200),
(42276),
(42351),
(42427),
(42502),
(42578),
(42654),
(42730),
(42806),
(42882),
(42959),
(43035),
(43111),
(43188),
(43265),
(43341),
(43418),
(43495),
(43572),
(43649),
(43727),
(43804),
(43882),
(43959),
(44037),
(44115),
(44192),
(44270),
(44349),
(44427),
(44505),
(44583),
(44662),
(44740),
(44819),
(44898),
(44977),
(45056),
(45135),
(45214),
(45293),
(45373),
(45452),
(45532),
(45612),
(45692),
(45771),
(45852),
(45932),
(46012),
(46092),
(46173),
(46253),
(46334),
(46415),
(46495),
(46576),
(46658),
(46739),
(46820),
(46901),
(46983),
(47064),
(47146),
(47228),
(47310),
(47392),
(47474),
(47556),
(47638),
(47721),
(47803),
(47886),
(47969),
(48052),
(48135),
(48218),
(48301),
(48384),
(48467),
(48551),
(48635),
(48718),
(48802),
(48886),
(48970),
(49054),
(49138),
(49223),
(49307),
(49392),
(49476),
(49561),
(49646),
(49731),
(49816),
(49901),
(49987),
(50072),
(50157),
(50243),
(50329),
(50415),
(50501),
(50587),
(50673),
(50759),
(50846),
(50932),
(51019),
(51105),
(51192),
(51279),
(51366),
(51453),
(51541),
(51628),
(51715),
(51803),
(51891),
(51978),
(52066),
(52154),
(52243),
(52331),
(52419),
(52508),
(52596),
(52685),
(52774),
(52863),
(52952),
(53041),
(53130),
(53219),
(53309),
(53398),
(53488),
(53578),
(53668),
(53758),
(53848),
(53938),
(54028),
(54119),
(54209),
(54300),
(54391),
(54482),
(54573),
(54664),
(54755),
(54847),
(54938),
(55030),
(55121),
(55213),
(55305),
(55397),
(55489),
(55582),
(55674),
(55766),
(55859),
(55952),
(56045),
(56138),
(56231),
(56324),
(56417),
(56510),
(56604),
(56698),
(56791),
(56885),
(56979),
(57073),
(57167),
(57262),
(57356),
(57451),
(57545),
(57640),
(57735),
(57830),
(57925),
(58021),
(58116),
(58211),
(58307),
(58403),
(58498),
(58594),
(58690),
(58787),
(58883),
(58979),
(59076),
(59173),
(59269),
(59366),
(59463),
(59560),
(59657),
(59755),
(59852),
(59950),
(60048),
(60145),
(60243),
(60341),
(60439),
(60538),
(60636),
(60735),
(60833),
(60932),
(61031),
(61130),
(61229),
(61328),
(61428),
(61527),
(61627),
(61726),
(61826),
(61926),
(62026),
(62126),
(62227),
(62327),
(62428),
(62528),
(62629),
(62730),
(62831),
(62932),
(63034),
(63135),
(63236),
(63338),
(63440),
(63542),
(63644),
(63746),
(63848),
(63950),
(64053),
(64155),
(64258),
(64361),
(64464),
(64567)  -- array index 4095 (voltage = "111111111111" or 4095 mV), distance output 3787 (37.87 cm)
);


end package LUT_pkg;
